module NV_NVDLA_CSC_WL_dec( // @[:@3.2]

  input          nvdla_core_clk, // @[:@6.4]
  input          nvdla_core_rstn, // @[:@6.4]
  input          input_pipe_valid, // @[:@6.4]
  input  [63:0]  input_mask, // @[:@6.4]
  input  [511:0] input_data, // @[:@6.4]
  input  [31:0]  input_sel, // @[:@6.4]
  input  [9:0]   input_mask_en, // @[:@6.4]
  output         output_pvld, // @[:@6.4]
  output [63:0]  output_mask, // @[:@6.4]
  output [7:0]   output_data0, // @[:@6.4]
  output [7:0]   output_data1, // @[:@6.4]
  output [7:0]   output_data2, // @[:@6.4]
  output [7:0]   output_data3, // @[:@6.4]
  output [7:0]   output_data4, // @[:@6.4]
  output [7:0]   output_data5, // @[:@6.4]
  output [7:0]   output_data6, // @[:@6.4]
  output [7:0]   output_data7, // @[:@6.4]
  output [7:0]   output_data8, // @[:@6.4]
  output [7:0]   output_data9, // @[:@6.4]
  output [7:0]   output_data10, // @[:@6.4]
  output [7:0]   output_data11, // @[:@6.4]
  output [7:0]   output_data12, // @[:@6.4]
  output [7:0]   output_data13, // @[:@6.4]
  output [7:0]   output_data14, // @[:@6.4]
  output [7:0]   output_data15, // @[:@6.4]
  output [7:0]   output_data16, // @[:@6.4]
  output [7:0]   output_data17, // @[:@6.4]
  output [7:0]   output_data18, // @[:@6.4]
  output [7:0]   output_data19, // @[:@6.4]
  output [7:0]   output_data20, // @[:@6.4]
  output [7:0]   output_data21, // @[:@6.4]
  output [7:0]   output_data22, // @[:@6.4]
  output [7:0]   output_data23, // @[:@6.4]
  output [7:0]   output_data24, // @[:@6.4]
  output [7:0]   output_data25, // @[:@6.4]
  output [7:0]   output_data26, // @[:@6.4]
  output [7:0]   output_data27, // @[:@6.4]
  output [7:0]   output_data28, // @[:@6.4]
  output [7:0]   output_data29, // @[:@6.4]
  output [7:0]   output_data30, // @[:@6.4]
  output [7:0]   output_data31, // @[:@6.4]
  output [7:0]   output_data32, // @[:@6.4]
  output [7:0]   output_data33, // @[:@6.4]
  output [7:0]   output_data34, // @[:@6.4]
  output [7:0]   output_data35, // @[:@6.4]
  output [7:0]   output_data36, // @[:@6.4]
  output [7:0]   output_data37, // @[:@6.4]
  output [7:0]   output_data38, // @[:@6.4]
  output [7:0]   output_data39, // @[:@6.4]
  output [7:0]   output_data40, // @[:@6.4]
  output [7:0]   output_data41, // @[:@6.4]
  output [7:0]   output_data42, // @[:@6.4]
  output [7:0]   output_data43, // @[:@6.4]
  output [7:0]   output_data44, // @[:@6.4]
  output [7:0]   output_data45, // @[:@6.4]
  output [7:0]   output_data46, // @[:@6.4]
  output [7:0]   output_data47, // @[:@6.4]
  output [7:0]   output_data48, // @[:@6.4]
  output [7:0]   output_data49, // @[:@6.4]
  output [7:0]   output_data50, // @[:@6.4]
  output [7:0]   output_data51, // @[:@6.4]
  output [7:0]   output_data52, // @[:@6.4]
  output [7:0]   output_data53, // @[:@6.4]
  output [7:0]   output_data54, // @[:@6.4]
  output [7:0]   output_data55, // @[:@6.4]
  output [7:0]   output_data56, // @[:@6.4]
  output [7:0]   output_data57, // @[:@6.4]
  output [7:0]   output_data58, // @[:@6.4]
  output [7:0]   output_data59, // @[:@6.4]
  output [7:0]   output_data60, // @[:@6.4]
  output [7:0]   output_data61, // @[:@6.4]
  output [7:0]   output_data62, // @[:@6.4]
  output [7:0]   output_data63, // @[:@6.4]
  output [31:0]  output_sel // @[:@6.4]
);
  wire  _T_326; // @[NV_NVDLA_CSC_WL_dec.scala 55:37:@8.4]
  wire  _T_397; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@10.4]
  wire  _T_398; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@12.4]
  wire  _T_399; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@14.4]
  wire  _T_400; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@16.4]
  wire  _T_401; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@18.4]
  wire  _T_402; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@20.4]
  wire  _T_403; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@22.4]
  wire  _T_404; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@24.4]
  wire  _T_405; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@26.4]
  wire  _T_406; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@28.4]
  wire  _T_407; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@30.4]
  wire  _T_408; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@32.4]
  wire  _T_409; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@34.4]
  wire  _T_410; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@36.4]
  wire  _T_411; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@38.4]
  wire  _T_412; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@40.4]
  wire  _T_413; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@42.4]
  wire  _T_414; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@44.4]
  wire  _T_415; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@46.4]
  wire  _T_416; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@48.4]
  wire  _T_417; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@50.4]
  wire  _T_418; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@52.4]
  wire  _T_419; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@54.4]
  wire  _T_420; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@56.4]
  wire  _T_421; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@58.4]
  wire  _T_422; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@60.4]
  wire  _T_423; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@62.4]
  wire  _T_424; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@64.4]
  wire  _T_425; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@66.4]
  wire  _T_426; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@68.4]
  wire  _T_427; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@70.4]
  wire  _T_428; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@72.4]
  wire  _T_429; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@74.4]
  wire  _T_430; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@76.4]
  wire  _T_431; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@78.4]
  wire  _T_432; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@80.4]
  wire  _T_433; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@82.4]
  wire  _T_434; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@84.4]
  wire  _T_435; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@86.4]
  wire  _T_436; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@88.4]
  wire  _T_437; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@90.4]
  wire  _T_438; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@92.4]
  wire  _T_439; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@94.4]
  wire  _T_440; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@96.4]
  wire  _T_441; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@98.4]
  wire  _T_442; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@100.4]
  wire  _T_443; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@102.4]
  wire  _T_444; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@104.4]
  wire  _T_445; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@106.4]
  wire  _T_446; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@108.4]
  wire  _T_447; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@110.4]
  wire  _T_448; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@112.4]
  wire  _T_449; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@114.4]
  wire  _T_450; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@116.4]
  wire  _T_451; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@118.4]
  wire  _T_452; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@120.4]
  wire  _T_453; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@122.4]
  wire  _T_454; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@124.4]
  wire  _T_455; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@126.4]
  wire  _T_456; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@128.4]
  wire  _T_457; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@130.4]
  wire  _T_458; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@132.4]
  wire  _T_459; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@134.4]
  wire  _T_460; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@136.4]
  wire [7:0] _T_531; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@139.4]
  wire [7:0] _T_532; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@141.4]
  wire [7:0] _T_533; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@143.4]
  wire [7:0] _T_534; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@145.4]
  wire [7:0] _T_535; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@147.4]
  wire [7:0] _T_536; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@149.4]
  wire [7:0] _T_537; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@151.4]
  wire [7:0] _T_538; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@153.4]
  wire [7:0] _T_539; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@155.4]
  wire [7:0] _T_540; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@157.4]
  wire [7:0] _T_541; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@159.4]
  wire [7:0] _T_542; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@161.4]
  wire [7:0] _T_543; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@163.4]
  wire [7:0] _T_544; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@165.4]
  wire [7:0] _T_545; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@167.4]
  wire [7:0] _T_546; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@169.4]
  wire [7:0] _T_547; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@171.4]
  wire [7:0] _T_548; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@173.4]
  wire [7:0] _T_549; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@175.4]
  wire [7:0] _T_550; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@177.4]
  wire [7:0] _T_551; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@179.4]
  wire [7:0] _T_552; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@181.4]
  wire [7:0] _T_553; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@183.4]
  wire [7:0] _T_554; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@185.4]
  wire [7:0] _T_555; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@187.4]
  wire [7:0] _T_556; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@189.4]
  wire [7:0] _T_557; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@191.4]
  wire [7:0] _T_558; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@193.4]
  wire [7:0] _T_559; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@195.4]
  wire [7:0] _T_560; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@197.4]
  wire [7:0] _T_561; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@199.4]
  wire [7:0] _T_562; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@201.4]
  wire [7:0] _T_563; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@203.4]
  wire [7:0] _T_564; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@205.4]
  wire [7:0] _T_565; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@207.4]
  wire [7:0] _T_566; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@209.4]
  wire [7:0] _T_567; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@211.4]
  wire [7:0] _T_568; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@213.4]
  wire [7:0] _T_569; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@215.4]
  wire [7:0] _T_570; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@217.4]
  wire [7:0] _T_571; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@219.4]
  wire [7:0] _T_572; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@221.4]
  wire [7:0] _T_573; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@223.4]
  wire [7:0] _T_574; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@225.4]
  wire [7:0] _T_575; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@227.4]
  wire [7:0] _T_576; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@229.4]
  wire [7:0] _T_577; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@231.4]
  wire [7:0] _T_578; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@233.4]
  wire [7:0] _T_579; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@235.4]
  wire [7:0] _T_580; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@237.4]
  wire [7:0] _T_581; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@239.4]
  wire [7:0] _T_582; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@241.4]
  wire [7:0] _T_583; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@243.4]
  wire [7:0] _T_584; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@245.4]
  wire [7:0] _T_585; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@247.4]
  wire [7:0] _T_586; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@249.4]
  wire [7:0] _T_587; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@251.4]
  wire [7:0] _T_588; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@253.4]
  wire [7:0] _T_589; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@255.4]
  wire [7:0] _T_590; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@257.4]
  wire [7:0] _T_591; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@259.4]
  wire [7:0] _T_592; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@261.4]
  wire [7:0] _T_593; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@263.4]
  wire [7:0] _T_594; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@265.4]
  wire  _T_633; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@268.4]
  wire  _T_634; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@270.4]
  wire  _T_635; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@272.4]
  wire  _T_636; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@274.4]
  wire  _T_637; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@276.4]
  wire  _T_638; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@278.4]
  wire  _T_639; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@280.4]
  wire  _T_640; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@282.4]
  wire  _T_641; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@284.4]
  wire  _T_642; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@286.4]
  wire  _T_643; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@288.4]
  wire  _T_644; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@290.4]
  wire  _T_645; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@292.4]
  wire  _T_646; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@294.4]
  wire  _T_647; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@296.4]
  wire  _T_648; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@298.4]
  wire  _T_649; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@300.4]
  wire  _T_650; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@302.4]
  wire  _T_651; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@304.4]
  wire  _T_652; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@306.4]
  wire  _T_653; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@308.4]
  wire  _T_654; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@310.4]
  wire  _T_655; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@312.4]
  wire  _T_656; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@314.4]
  wire  _T_657; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@316.4]
  wire  _T_658; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@318.4]
  wire  _T_659; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@320.4]
  wire  _T_660; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@322.4]
  wire  _T_661; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@324.4]
  wire  _T_662; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@326.4]
  wire  _T_663; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@328.4]
  wire  _T_664; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@330.4]
  wire  _T_665; // @[NV_NVDLA_CSC_WL_dec.scala 81:48:@332.4]
  wire  _T_800_0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_1; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_2; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_3; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_4; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_5; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_6; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_7; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_8; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_9; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_10; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_11; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_12; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_13; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_14; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_15; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_16; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_17; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_18; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_19; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_20; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_21; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_22; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_23; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_24; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_25; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_26; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_27; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_28; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_29; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_30; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_31; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_32; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_33; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_34; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_35; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_36; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_37; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_38; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_39; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_40; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_41; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_42; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_43; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_44; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_45; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_46; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_47; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_48; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_49; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_50; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_51; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_52; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_53; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_54; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_55; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_56; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_57; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_58; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_59; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_60; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_61; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_62; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire  _T_800_63; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  wire [7:0] _T_1068; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@406.4]
  wire [15:0] _T_1076; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@414.4]
  wire [7:0] _T_1083; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@421.4]
  wire [31:0] _T_1092; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@430.4]
  wire [7:0] _T_1099; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@437.4]
  wire [15:0] _T_1107; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@445.4]
  wire [7:0] _T_1114; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@452.4]
  wire [31:0] _T_1123; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@461.4]
  wire [63:0] _T_1124; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@462.4]
  wire  _T_1125; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@463.4]
  wire [1:0] _T_1190; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@529.4]
  wire  _T_1191; // @[Bitwise.scala 50:65:@530.4]
  wire  _T_1192; // @[Bitwise.scala 50:65:@531.4]
  wire [1:0] _T_1193; // @[Bitwise.scala 48:55:@532.4]
  wire [2:0] _T_1257; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@597.4]
  wire  _T_1258; // @[Bitwise.scala 50:65:@598.4]
  wire  _T_1259; // @[Bitwise.scala 50:65:@599.4]
  wire  _T_1260; // @[Bitwise.scala 50:65:@600.4]
  wire [1:0] _T_1261; // @[Bitwise.scala 48:55:@601.4]
  wire [1:0] _GEN_544; // @[Bitwise.scala 48:55:@602.4]
  wire [2:0] _T_1262; // @[Bitwise.scala 48:55:@602.4]
  wire [3:0] _T_1326; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@667.4]
  wire  _T_1327; // @[Bitwise.scala 50:65:@668.4]
  wire  _T_1328; // @[Bitwise.scala 50:65:@669.4]
  wire  _T_1329; // @[Bitwise.scala 50:65:@670.4]
  wire  _T_1330; // @[Bitwise.scala 50:65:@671.4]
  wire [1:0] _T_1331; // @[Bitwise.scala 48:55:@672.4]
  wire [1:0] _T_1332; // @[Bitwise.scala 48:55:@673.4]
  wire [2:0] _T_1333; // @[Bitwise.scala 48:55:@674.4]
  wire [4:0] _T_1397; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@739.4]
  wire  _T_1398; // @[Bitwise.scala 50:65:@740.4]
  wire  _T_1399; // @[Bitwise.scala 50:65:@741.4]
  wire  _T_1400; // @[Bitwise.scala 50:65:@742.4]
  wire  _T_1401; // @[Bitwise.scala 50:65:@743.4]
  wire  _T_1402; // @[Bitwise.scala 50:65:@744.4]
  wire [1:0] _T_1403; // @[Bitwise.scala 48:55:@745.4]
  wire [1:0] _T_1404; // @[Bitwise.scala 48:55:@746.4]
  wire [1:0] _GEN_545; // @[Bitwise.scala 48:55:@747.4]
  wire [2:0] _T_1405; // @[Bitwise.scala 48:55:@747.4]
  wire [2:0] _GEN_546; // @[Bitwise.scala 48:55:@748.4]
  wire [3:0] _T_1406; // @[Bitwise.scala 48:55:@748.4]
  wire [5:0] _T_1470; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@813.4]
  wire  _T_1471; // @[Bitwise.scala 50:65:@814.4]
  wire  _T_1472; // @[Bitwise.scala 50:65:@815.4]
  wire  _T_1473; // @[Bitwise.scala 50:65:@816.4]
  wire  _T_1474; // @[Bitwise.scala 50:65:@817.4]
  wire  _T_1475; // @[Bitwise.scala 50:65:@818.4]
  wire  _T_1476; // @[Bitwise.scala 50:65:@819.4]
  wire [1:0] _T_1477; // @[Bitwise.scala 48:55:@820.4]
  wire [1:0] _GEN_547; // @[Bitwise.scala 48:55:@821.4]
  wire [2:0] _T_1478; // @[Bitwise.scala 48:55:@821.4]
  wire [1:0] _T_1479; // @[Bitwise.scala 48:55:@822.4]
  wire [1:0] _GEN_548; // @[Bitwise.scala 48:55:@823.4]
  wire [2:0] _T_1480; // @[Bitwise.scala 48:55:@823.4]
  wire [3:0] _T_1481; // @[Bitwise.scala 48:55:@824.4]
  wire [6:0] _T_1545; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@889.4]
  wire  _T_1546; // @[Bitwise.scala 50:65:@890.4]
  wire  _T_1547; // @[Bitwise.scala 50:65:@891.4]
  wire  _T_1548; // @[Bitwise.scala 50:65:@892.4]
  wire  _T_1549; // @[Bitwise.scala 50:65:@893.4]
  wire  _T_1550; // @[Bitwise.scala 50:65:@894.4]
  wire  _T_1551; // @[Bitwise.scala 50:65:@895.4]
  wire  _T_1552; // @[Bitwise.scala 50:65:@896.4]
  wire [1:0] _T_1553; // @[Bitwise.scala 48:55:@897.4]
  wire [1:0] _GEN_549; // @[Bitwise.scala 48:55:@898.4]
  wire [2:0] _T_1554; // @[Bitwise.scala 48:55:@898.4]
  wire [1:0] _T_1555; // @[Bitwise.scala 48:55:@899.4]
  wire [1:0] _T_1556; // @[Bitwise.scala 48:55:@900.4]
  wire [2:0] _T_1557; // @[Bitwise.scala 48:55:@901.4]
  wire [3:0] _T_1558; // @[Bitwise.scala 48:55:@902.4]
  wire [7:0] _T_1622; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@967.4]
  wire  _T_1623; // @[Bitwise.scala 50:65:@968.4]
  wire  _T_1624; // @[Bitwise.scala 50:65:@969.4]
  wire  _T_1625; // @[Bitwise.scala 50:65:@970.4]
  wire  _T_1626; // @[Bitwise.scala 50:65:@971.4]
  wire  _T_1627; // @[Bitwise.scala 50:65:@972.4]
  wire  _T_1628; // @[Bitwise.scala 50:65:@973.4]
  wire  _T_1629; // @[Bitwise.scala 50:65:@974.4]
  wire  _T_1630; // @[Bitwise.scala 50:65:@975.4]
  wire [1:0] _T_1631; // @[Bitwise.scala 48:55:@976.4]
  wire [1:0] _T_1632; // @[Bitwise.scala 48:55:@977.4]
  wire [2:0] _T_1633; // @[Bitwise.scala 48:55:@978.4]
  wire [1:0] _T_1634; // @[Bitwise.scala 48:55:@979.4]
  wire [1:0] _T_1635; // @[Bitwise.scala 48:55:@980.4]
  wire [2:0] _T_1636; // @[Bitwise.scala 48:55:@981.4]
  wire [3:0] _T_1637; // @[Bitwise.scala 48:55:@982.4]
  wire [8:0] _T_1701; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1047.4]
  wire  _T_1702; // @[Bitwise.scala 50:65:@1048.4]
  wire  _T_1703; // @[Bitwise.scala 50:65:@1049.4]
  wire  _T_1704; // @[Bitwise.scala 50:65:@1050.4]
  wire  _T_1705; // @[Bitwise.scala 50:65:@1051.4]
  wire  _T_1706; // @[Bitwise.scala 50:65:@1052.4]
  wire  _T_1707; // @[Bitwise.scala 50:65:@1053.4]
  wire  _T_1708; // @[Bitwise.scala 50:65:@1054.4]
  wire  _T_1709; // @[Bitwise.scala 50:65:@1055.4]
  wire  _T_1710; // @[Bitwise.scala 50:65:@1056.4]
  wire [1:0] _T_1711; // @[Bitwise.scala 48:55:@1057.4]
  wire [1:0] _T_1712; // @[Bitwise.scala 48:55:@1058.4]
  wire [2:0] _T_1713; // @[Bitwise.scala 48:55:@1059.4]
  wire [1:0] _T_1714; // @[Bitwise.scala 48:55:@1060.4]
  wire [1:0] _T_1715; // @[Bitwise.scala 48:55:@1061.4]
  wire [1:0] _GEN_550; // @[Bitwise.scala 48:55:@1062.4]
  wire [2:0] _T_1716; // @[Bitwise.scala 48:55:@1062.4]
  wire [2:0] _GEN_551; // @[Bitwise.scala 48:55:@1063.4]
  wire [3:0] _T_1717; // @[Bitwise.scala 48:55:@1063.4]
  wire [3:0] _GEN_552; // @[Bitwise.scala 48:55:@1064.4]
  wire [4:0] _T_1718; // @[Bitwise.scala 48:55:@1064.4]
  wire [9:0] _T_1782; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1129.4]
  wire  _T_1783; // @[Bitwise.scala 50:65:@1130.4]
  wire  _T_1784; // @[Bitwise.scala 50:65:@1131.4]
  wire  _T_1785; // @[Bitwise.scala 50:65:@1132.4]
  wire  _T_1786; // @[Bitwise.scala 50:65:@1133.4]
  wire  _T_1787; // @[Bitwise.scala 50:65:@1134.4]
  wire  _T_1788; // @[Bitwise.scala 50:65:@1135.4]
  wire  _T_1789; // @[Bitwise.scala 50:65:@1136.4]
  wire  _T_1790; // @[Bitwise.scala 50:65:@1137.4]
  wire  _T_1791; // @[Bitwise.scala 50:65:@1138.4]
  wire  _T_1792; // @[Bitwise.scala 50:65:@1139.4]
  wire [1:0] _T_1793; // @[Bitwise.scala 48:55:@1140.4]
  wire [1:0] _T_1794; // @[Bitwise.scala 48:55:@1141.4]
  wire [1:0] _GEN_553; // @[Bitwise.scala 48:55:@1142.4]
  wire [2:0] _T_1795; // @[Bitwise.scala 48:55:@1142.4]
  wire [2:0] _GEN_554; // @[Bitwise.scala 48:55:@1143.4]
  wire [3:0] _T_1796; // @[Bitwise.scala 48:55:@1143.4]
  wire [1:0] _T_1797; // @[Bitwise.scala 48:55:@1144.4]
  wire [1:0] _T_1798; // @[Bitwise.scala 48:55:@1145.4]
  wire [1:0] _GEN_555; // @[Bitwise.scala 48:55:@1146.4]
  wire [2:0] _T_1799; // @[Bitwise.scala 48:55:@1146.4]
  wire [2:0] _GEN_556; // @[Bitwise.scala 48:55:@1147.4]
  wire [3:0] _T_1800; // @[Bitwise.scala 48:55:@1147.4]
  wire [4:0] _T_1801; // @[Bitwise.scala 48:55:@1148.4]
  wire [10:0] _T_1865; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1213.4]
  wire  _T_1866; // @[Bitwise.scala 50:65:@1214.4]
  wire  _T_1867; // @[Bitwise.scala 50:65:@1215.4]
  wire  _T_1868; // @[Bitwise.scala 50:65:@1216.4]
  wire  _T_1869; // @[Bitwise.scala 50:65:@1217.4]
  wire  _T_1870; // @[Bitwise.scala 50:65:@1218.4]
  wire  _T_1871; // @[Bitwise.scala 50:65:@1219.4]
  wire  _T_1872; // @[Bitwise.scala 50:65:@1220.4]
  wire  _T_1873; // @[Bitwise.scala 50:65:@1221.4]
  wire  _T_1874; // @[Bitwise.scala 50:65:@1222.4]
  wire  _T_1875; // @[Bitwise.scala 50:65:@1223.4]
  wire  _T_1876; // @[Bitwise.scala 50:65:@1224.4]
  wire [1:0] _T_1877; // @[Bitwise.scala 48:55:@1225.4]
  wire [1:0] _T_1878; // @[Bitwise.scala 48:55:@1226.4]
  wire [1:0] _GEN_557; // @[Bitwise.scala 48:55:@1227.4]
  wire [2:0] _T_1879; // @[Bitwise.scala 48:55:@1227.4]
  wire [2:0] _GEN_558; // @[Bitwise.scala 48:55:@1228.4]
  wire [3:0] _T_1880; // @[Bitwise.scala 48:55:@1228.4]
  wire [1:0] _T_1881; // @[Bitwise.scala 48:55:@1229.4]
  wire [1:0] _GEN_559; // @[Bitwise.scala 48:55:@1230.4]
  wire [2:0] _T_1882; // @[Bitwise.scala 48:55:@1230.4]
  wire [1:0] _T_1883; // @[Bitwise.scala 48:55:@1231.4]
  wire [1:0] _GEN_560; // @[Bitwise.scala 48:55:@1232.4]
  wire [2:0] _T_1884; // @[Bitwise.scala 48:55:@1232.4]
  wire [3:0] _T_1885; // @[Bitwise.scala 48:55:@1233.4]
  wire [4:0] _T_1886; // @[Bitwise.scala 48:55:@1234.4]
  wire [11:0] _T_1950; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1299.4]
  wire  _T_1951; // @[Bitwise.scala 50:65:@1300.4]
  wire  _T_1952; // @[Bitwise.scala 50:65:@1301.4]
  wire  _T_1953; // @[Bitwise.scala 50:65:@1302.4]
  wire  _T_1954; // @[Bitwise.scala 50:65:@1303.4]
  wire  _T_1955; // @[Bitwise.scala 50:65:@1304.4]
  wire  _T_1956; // @[Bitwise.scala 50:65:@1305.4]
  wire  _T_1957; // @[Bitwise.scala 50:65:@1306.4]
  wire  _T_1958; // @[Bitwise.scala 50:65:@1307.4]
  wire  _T_1959; // @[Bitwise.scala 50:65:@1308.4]
  wire  _T_1960; // @[Bitwise.scala 50:65:@1309.4]
  wire  _T_1961; // @[Bitwise.scala 50:65:@1310.4]
  wire  _T_1962; // @[Bitwise.scala 50:65:@1311.4]
  wire [1:0] _T_1963; // @[Bitwise.scala 48:55:@1312.4]
  wire [1:0] _GEN_561; // @[Bitwise.scala 48:55:@1313.4]
  wire [2:0] _T_1964; // @[Bitwise.scala 48:55:@1313.4]
  wire [1:0] _T_1965; // @[Bitwise.scala 48:55:@1314.4]
  wire [1:0] _GEN_562; // @[Bitwise.scala 48:55:@1315.4]
  wire [2:0] _T_1966; // @[Bitwise.scala 48:55:@1315.4]
  wire [3:0] _T_1967; // @[Bitwise.scala 48:55:@1316.4]
  wire [1:0] _T_1968; // @[Bitwise.scala 48:55:@1317.4]
  wire [1:0] _GEN_563; // @[Bitwise.scala 48:55:@1318.4]
  wire [2:0] _T_1969; // @[Bitwise.scala 48:55:@1318.4]
  wire [1:0] _T_1970; // @[Bitwise.scala 48:55:@1319.4]
  wire [1:0] _GEN_564; // @[Bitwise.scala 48:55:@1320.4]
  wire [2:0] _T_1971; // @[Bitwise.scala 48:55:@1320.4]
  wire [3:0] _T_1972; // @[Bitwise.scala 48:55:@1321.4]
  wire [4:0] _T_1973; // @[Bitwise.scala 48:55:@1322.4]
  wire [12:0] _T_2037; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1387.4]
  wire  _T_2038; // @[Bitwise.scala 50:65:@1388.4]
  wire  _T_2039; // @[Bitwise.scala 50:65:@1389.4]
  wire  _T_2040; // @[Bitwise.scala 50:65:@1390.4]
  wire  _T_2041; // @[Bitwise.scala 50:65:@1391.4]
  wire  _T_2042; // @[Bitwise.scala 50:65:@1392.4]
  wire  _T_2043; // @[Bitwise.scala 50:65:@1393.4]
  wire  _T_2044; // @[Bitwise.scala 50:65:@1394.4]
  wire  _T_2045; // @[Bitwise.scala 50:65:@1395.4]
  wire  _T_2046; // @[Bitwise.scala 50:65:@1396.4]
  wire  _T_2047; // @[Bitwise.scala 50:65:@1397.4]
  wire  _T_2048; // @[Bitwise.scala 50:65:@1398.4]
  wire  _T_2049; // @[Bitwise.scala 50:65:@1399.4]
  wire  _T_2050; // @[Bitwise.scala 50:65:@1400.4]
  wire [1:0] _T_2051; // @[Bitwise.scala 48:55:@1401.4]
  wire [1:0] _GEN_565; // @[Bitwise.scala 48:55:@1402.4]
  wire [2:0] _T_2052; // @[Bitwise.scala 48:55:@1402.4]
  wire [1:0] _T_2053; // @[Bitwise.scala 48:55:@1403.4]
  wire [1:0] _GEN_566; // @[Bitwise.scala 48:55:@1404.4]
  wire [2:0] _T_2054; // @[Bitwise.scala 48:55:@1404.4]
  wire [3:0] _T_2055; // @[Bitwise.scala 48:55:@1405.4]
  wire [1:0] _T_2056; // @[Bitwise.scala 48:55:@1406.4]
  wire [1:0] _GEN_567; // @[Bitwise.scala 48:55:@1407.4]
  wire [2:0] _T_2057; // @[Bitwise.scala 48:55:@1407.4]
  wire [1:0] _T_2058; // @[Bitwise.scala 48:55:@1408.4]
  wire [1:0] _T_2059; // @[Bitwise.scala 48:55:@1409.4]
  wire [2:0] _T_2060; // @[Bitwise.scala 48:55:@1410.4]
  wire [3:0] _T_2061; // @[Bitwise.scala 48:55:@1411.4]
  wire [4:0] _T_2062; // @[Bitwise.scala 48:55:@1412.4]
  wire [13:0] _T_2126; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1477.4]
  wire  _T_2127; // @[Bitwise.scala 50:65:@1478.4]
  wire  _T_2128; // @[Bitwise.scala 50:65:@1479.4]
  wire  _T_2129; // @[Bitwise.scala 50:65:@1480.4]
  wire  _T_2130; // @[Bitwise.scala 50:65:@1481.4]
  wire  _T_2131; // @[Bitwise.scala 50:65:@1482.4]
  wire  _T_2132; // @[Bitwise.scala 50:65:@1483.4]
  wire  _T_2133; // @[Bitwise.scala 50:65:@1484.4]
  wire  _T_2134; // @[Bitwise.scala 50:65:@1485.4]
  wire  _T_2135; // @[Bitwise.scala 50:65:@1486.4]
  wire  _T_2136; // @[Bitwise.scala 50:65:@1487.4]
  wire  _T_2137; // @[Bitwise.scala 50:65:@1488.4]
  wire  _T_2138; // @[Bitwise.scala 50:65:@1489.4]
  wire  _T_2139; // @[Bitwise.scala 50:65:@1490.4]
  wire  _T_2140; // @[Bitwise.scala 50:65:@1491.4]
  wire [1:0] _T_2141; // @[Bitwise.scala 48:55:@1492.4]
  wire [1:0] _GEN_568; // @[Bitwise.scala 48:55:@1493.4]
  wire [2:0] _T_2142; // @[Bitwise.scala 48:55:@1493.4]
  wire [1:0] _T_2143; // @[Bitwise.scala 48:55:@1494.4]
  wire [1:0] _T_2144; // @[Bitwise.scala 48:55:@1495.4]
  wire [2:0] _T_2145; // @[Bitwise.scala 48:55:@1496.4]
  wire [3:0] _T_2146; // @[Bitwise.scala 48:55:@1497.4]
  wire [1:0] _T_2147; // @[Bitwise.scala 48:55:@1498.4]
  wire [1:0] _GEN_569; // @[Bitwise.scala 48:55:@1499.4]
  wire [2:0] _T_2148; // @[Bitwise.scala 48:55:@1499.4]
  wire [1:0] _T_2149; // @[Bitwise.scala 48:55:@1500.4]
  wire [1:0] _T_2150; // @[Bitwise.scala 48:55:@1501.4]
  wire [2:0] _T_2151; // @[Bitwise.scala 48:55:@1502.4]
  wire [3:0] _T_2152; // @[Bitwise.scala 48:55:@1503.4]
  wire [4:0] _T_2153; // @[Bitwise.scala 48:55:@1504.4]
  wire [14:0] _T_2217; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1569.4]
  wire  _T_2218; // @[Bitwise.scala 50:65:@1570.4]
  wire  _T_2219; // @[Bitwise.scala 50:65:@1571.4]
  wire  _T_2220; // @[Bitwise.scala 50:65:@1572.4]
  wire  _T_2221; // @[Bitwise.scala 50:65:@1573.4]
  wire  _T_2222; // @[Bitwise.scala 50:65:@1574.4]
  wire  _T_2223; // @[Bitwise.scala 50:65:@1575.4]
  wire  _T_2224; // @[Bitwise.scala 50:65:@1576.4]
  wire  _T_2225; // @[Bitwise.scala 50:65:@1577.4]
  wire  _T_2226; // @[Bitwise.scala 50:65:@1578.4]
  wire  _T_2227; // @[Bitwise.scala 50:65:@1579.4]
  wire  _T_2228; // @[Bitwise.scala 50:65:@1580.4]
  wire  _T_2229; // @[Bitwise.scala 50:65:@1581.4]
  wire  _T_2230; // @[Bitwise.scala 50:65:@1582.4]
  wire  _T_2231; // @[Bitwise.scala 50:65:@1583.4]
  wire  _T_2232; // @[Bitwise.scala 50:65:@1584.4]
  wire [1:0] _T_2233; // @[Bitwise.scala 48:55:@1585.4]
  wire [1:0] _GEN_570; // @[Bitwise.scala 48:55:@1586.4]
  wire [2:0] _T_2234; // @[Bitwise.scala 48:55:@1586.4]
  wire [1:0] _T_2235; // @[Bitwise.scala 48:55:@1587.4]
  wire [1:0] _T_2236; // @[Bitwise.scala 48:55:@1588.4]
  wire [2:0] _T_2237; // @[Bitwise.scala 48:55:@1589.4]
  wire [3:0] _T_2238; // @[Bitwise.scala 48:55:@1590.4]
  wire [1:0] _T_2239; // @[Bitwise.scala 48:55:@1591.4]
  wire [1:0] _T_2240; // @[Bitwise.scala 48:55:@1592.4]
  wire [2:0] _T_2241; // @[Bitwise.scala 48:55:@1593.4]
  wire [1:0] _T_2242; // @[Bitwise.scala 48:55:@1594.4]
  wire [1:0] _T_2243; // @[Bitwise.scala 48:55:@1595.4]
  wire [2:0] _T_2244; // @[Bitwise.scala 48:55:@1596.4]
  wire [3:0] _T_2245; // @[Bitwise.scala 48:55:@1597.4]
  wire [4:0] _T_2246; // @[Bitwise.scala 48:55:@1598.4]
  wire [15:0] _T_2310; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1663.4]
  wire  _T_2311; // @[Bitwise.scala 50:65:@1664.4]
  wire  _T_2312; // @[Bitwise.scala 50:65:@1665.4]
  wire  _T_2313; // @[Bitwise.scala 50:65:@1666.4]
  wire  _T_2314; // @[Bitwise.scala 50:65:@1667.4]
  wire  _T_2315; // @[Bitwise.scala 50:65:@1668.4]
  wire  _T_2316; // @[Bitwise.scala 50:65:@1669.4]
  wire  _T_2317; // @[Bitwise.scala 50:65:@1670.4]
  wire  _T_2318; // @[Bitwise.scala 50:65:@1671.4]
  wire  _T_2319; // @[Bitwise.scala 50:65:@1672.4]
  wire  _T_2320; // @[Bitwise.scala 50:65:@1673.4]
  wire  _T_2321; // @[Bitwise.scala 50:65:@1674.4]
  wire  _T_2322; // @[Bitwise.scala 50:65:@1675.4]
  wire  _T_2323; // @[Bitwise.scala 50:65:@1676.4]
  wire  _T_2324; // @[Bitwise.scala 50:65:@1677.4]
  wire  _T_2325; // @[Bitwise.scala 50:65:@1678.4]
  wire  _T_2326; // @[Bitwise.scala 50:65:@1679.4]
  wire [1:0] _T_2327; // @[Bitwise.scala 48:55:@1680.4]
  wire [1:0] _T_2328; // @[Bitwise.scala 48:55:@1681.4]
  wire [2:0] _T_2329; // @[Bitwise.scala 48:55:@1682.4]
  wire [1:0] _T_2330; // @[Bitwise.scala 48:55:@1683.4]
  wire [1:0] _T_2331; // @[Bitwise.scala 48:55:@1684.4]
  wire [2:0] _T_2332; // @[Bitwise.scala 48:55:@1685.4]
  wire [3:0] _T_2333; // @[Bitwise.scala 48:55:@1686.4]
  wire [1:0] _T_2334; // @[Bitwise.scala 48:55:@1687.4]
  wire [1:0] _T_2335; // @[Bitwise.scala 48:55:@1688.4]
  wire [2:0] _T_2336; // @[Bitwise.scala 48:55:@1689.4]
  wire [1:0] _T_2337; // @[Bitwise.scala 48:55:@1690.4]
  wire [1:0] _T_2338; // @[Bitwise.scala 48:55:@1691.4]
  wire [2:0] _T_2339; // @[Bitwise.scala 48:55:@1692.4]
  wire [3:0] _T_2340; // @[Bitwise.scala 48:55:@1693.4]
  wire [4:0] _T_2341; // @[Bitwise.scala 48:55:@1694.4]
  wire [16:0] _T_2405; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1759.4]
  wire  _T_2406; // @[Bitwise.scala 50:65:@1760.4]
  wire  _T_2407; // @[Bitwise.scala 50:65:@1761.4]
  wire  _T_2408; // @[Bitwise.scala 50:65:@1762.4]
  wire  _T_2409; // @[Bitwise.scala 50:65:@1763.4]
  wire  _T_2410; // @[Bitwise.scala 50:65:@1764.4]
  wire  _T_2411; // @[Bitwise.scala 50:65:@1765.4]
  wire  _T_2412; // @[Bitwise.scala 50:65:@1766.4]
  wire  _T_2413; // @[Bitwise.scala 50:65:@1767.4]
  wire  _T_2414; // @[Bitwise.scala 50:65:@1768.4]
  wire  _T_2415; // @[Bitwise.scala 50:65:@1769.4]
  wire  _T_2416; // @[Bitwise.scala 50:65:@1770.4]
  wire  _T_2417; // @[Bitwise.scala 50:65:@1771.4]
  wire  _T_2418; // @[Bitwise.scala 50:65:@1772.4]
  wire  _T_2419; // @[Bitwise.scala 50:65:@1773.4]
  wire  _T_2420; // @[Bitwise.scala 50:65:@1774.4]
  wire  _T_2421; // @[Bitwise.scala 50:65:@1775.4]
  wire  _T_2422; // @[Bitwise.scala 50:65:@1776.4]
  wire [1:0] _T_2423; // @[Bitwise.scala 48:55:@1777.4]
  wire [1:0] _T_2424; // @[Bitwise.scala 48:55:@1778.4]
  wire [2:0] _T_2425; // @[Bitwise.scala 48:55:@1779.4]
  wire [1:0] _T_2426; // @[Bitwise.scala 48:55:@1780.4]
  wire [1:0] _T_2427; // @[Bitwise.scala 48:55:@1781.4]
  wire [2:0] _T_2428; // @[Bitwise.scala 48:55:@1782.4]
  wire [3:0] _T_2429; // @[Bitwise.scala 48:55:@1783.4]
  wire [1:0] _T_2430; // @[Bitwise.scala 48:55:@1784.4]
  wire [1:0] _T_2431; // @[Bitwise.scala 48:55:@1785.4]
  wire [2:0] _T_2432; // @[Bitwise.scala 48:55:@1786.4]
  wire [1:0] _T_2433; // @[Bitwise.scala 48:55:@1787.4]
  wire [1:0] _T_2434; // @[Bitwise.scala 48:55:@1788.4]
  wire [1:0] _GEN_571; // @[Bitwise.scala 48:55:@1789.4]
  wire [2:0] _T_2435; // @[Bitwise.scala 48:55:@1789.4]
  wire [2:0] _GEN_572; // @[Bitwise.scala 48:55:@1790.4]
  wire [3:0] _T_2436; // @[Bitwise.scala 48:55:@1790.4]
  wire [3:0] _GEN_573; // @[Bitwise.scala 48:55:@1791.4]
  wire [4:0] _T_2437; // @[Bitwise.scala 48:55:@1791.4]
  wire [4:0] _GEN_574; // @[Bitwise.scala 48:55:@1792.4]
  wire [5:0] _T_2438; // @[Bitwise.scala 48:55:@1792.4]
  wire [17:0] _T_2502; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1857.4]
  wire  _T_2503; // @[Bitwise.scala 50:65:@1858.4]
  wire  _T_2504; // @[Bitwise.scala 50:65:@1859.4]
  wire  _T_2505; // @[Bitwise.scala 50:65:@1860.4]
  wire  _T_2506; // @[Bitwise.scala 50:65:@1861.4]
  wire  _T_2507; // @[Bitwise.scala 50:65:@1862.4]
  wire  _T_2508; // @[Bitwise.scala 50:65:@1863.4]
  wire  _T_2509; // @[Bitwise.scala 50:65:@1864.4]
  wire  _T_2510; // @[Bitwise.scala 50:65:@1865.4]
  wire  _T_2511; // @[Bitwise.scala 50:65:@1866.4]
  wire  _T_2512; // @[Bitwise.scala 50:65:@1867.4]
  wire  _T_2513; // @[Bitwise.scala 50:65:@1868.4]
  wire  _T_2514; // @[Bitwise.scala 50:65:@1869.4]
  wire  _T_2515; // @[Bitwise.scala 50:65:@1870.4]
  wire  _T_2516; // @[Bitwise.scala 50:65:@1871.4]
  wire  _T_2517; // @[Bitwise.scala 50:65:@1872.4]
  wire  _T_2518; // @[Bitwise.scala 50:65:@1873.4]
  wire  _T_2519; // @[Bitwise.scala 50:65:@1874.4]
  wire  _T_2520; // @[Bitwise.scala 50:65:@1875.4]
  wire [1:0] _T_2521; // @[Bitwise.scala 48:55:@1876.4]
  wire [1:0] _T_2522; // @[Bitwise.scala 48:55:@1877.4]
  wire [2:0] _T_2523; // @[Bitwise.scala 48:55:@1878.4]
  wire [1:0] _T_2524; // @[Bitwise.scala 48:55:@1879.4]
  wire [1:0] _T_2525; // @[Bitwise.scala 48:55:@1880.4]
  wire [1:0] _GEN_575; // @[Bitwise.scala 48:55:@1881.4]
  wire [2:0] _T_2526; // @[Bitwise.scala 48:55:@1881.4]
  wire [2:0] _GEN_576; // @[Bitwise.scala 48:55:@1882.4]
  wire [3:0] _T_2527; // @[Bitwise.scala 48:55:@1882.4]
  wire [3:0] _GEN_577; // @[Bitwise.scala 48:55:@1883.4]
  wire [4:0] _T_2528; // @[Bitwise.scala 48:55:@1883.4]
  wire [1:0] _T_2529; // @[Bitwise.scala 48:55:@1884.4]
  wire [1:0] _T_2530; // @[Bitwise.scala 48:55:@1885.4]
  wire [2:0] _T_2531; // @[Bitwise.scala 48:55:@1886.4]
  wire [1:0] _T_2532; // @[Bitwise.scala 48:55:@1887.4]
  wire [1:0] _T_2533; // @[Bitwise.scala 48:55:@1888.4]
  wire [1:0] _GEN_578; // @[Bitwise.scala 48:55:@1889.4]
  wire [2:0] _T_2534; // @[Bitwise.scala 48:55:@1889.4]
  wire [2:0] _GEN_579; // @[Bitwise.scala 48:55:@1890.4]
  wire [3:0] _T_2535; // @[Bitwise.scala 48:55:@1890.4]
  wire [3:0] _GEN_580; // @[Bitwise.scala 48:55:@1891.4]
  wire [4:0] _T_2536; // @[Bitwise.scala 48:55:@1891.4]
  wire [5:0] _T_2537; // @[Bitwise.scala 48:55:@1892.4]
  wire [18:0] _T_2601; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1957.4]
  wire  _T_2602; // @[Bitwise.scala 50:65:@1958.4]
  wire  _T_2603; // @[Bitwise.scala 50:65:@1959.4]
  wire  _T_2604; // @[Bitwise.scala 50:65:@1960.4]
  wire  _T_2605; // @[Bitwise.scala 50:65:@1961.4]
  wire  _T_2606; // @[Bitwise.scala 50:65:@1962.4]
  wire  _T_2607; // @[Bitwise.scala 50:65:@1963.4]
  wire  _T_2608; // @[Bitwise.scala 50:65:@1964.4]
  wire  _T_2609; // @[Bitwise.scala 50:65:@1965.4]
  wire  _T_2610; // @[Bitwise.scala 50:65:@1966.4]
  wire  _T_2611; // @[Bitwise.scala 50:65:@1967.4]
  wire  _T_2612; // @[Bitwise.scala 50:65:@1968.4]
  wire  _T_2613; // @[Bitwise.scala 50:65:@1969.4]
  wire  _T_2614; // @[Bitwise.scala 50:65:@1970.4]
  wire  _T_2615; // @[Bitwise.scala 50:65:@1971.4]
  wire  _T_2616; // @[Bitwise.scala 50:65:@1972.4]
  wire  _T_2617; // @[Bitwise.scala 50:65:@1973.4]
  wire  _T_2618; // @[Bitwise.scala 50:65:@1974.4]
  wire  _T_2619; // @[Bitwise.scala 50:65:@1975.4]
  wire  _T_2620; // @[Bitwise.scala 50:65:@1976.4]
  wire [1:0] _T_2621; // @[Bitwise.scala 48:55:@1977.4]
  wire [1:0] _T_2622; // @[Bitwise.scala 48:55:@1978.4]
  wire [2:0] _T_2623; // @[Bitwise.scala 48:55:@1979.4]
  wire [1:0] _T_2624; // @[Bitwise.scala 48:55:@1980.4]
  wire [1:0] _T_2625; // @[Bitwise.scala 48:55:@1981.4]
  wire [1:0] _GEN_581; // @[Bitwise.scala 48:55:@1982.4]
  wire [2:0] _T_2626; // @[Bitwise.scala 48:55:@1982.4]
  wire [2:0] _GEN_582; // @[Bitwise.scala 48:55:@1983.4]
  wire [3:0] _T_2627; // @[Bitwise.scala 48:55:@1983.4]
  wire [3:0] _GEN_583; // @[Bitwise.scala 48:55:@1984.4]
  wire [4:0] _T_2628; // @[Bitwise.scala 48:55:@1984.4]
  wire [1:0] _T_2629; // @[Bitwise.scala 48:55:@1985.4]
  wire [1:0] _T_2630; // @[Bitwise.scala 48:55:@1986.4]
  wire [1:0] _GEN_584; // @[Bitwise.scala 48:55:@1987.4]
  wire [2:0] _T_2631; // @[Bitwise.scala 48:55:@1987.4]
  wire [2:0] _GEN_585; // @[Bitwise.scala 48:55:@1988.4]
  wire [3:0] _T_2632; // @[Bitwise.scala 48:55:@1988.4]
  wire [1:0] _T_2633; // @[Bitwise.scala 48:55:@1989.4]
  wire [1:0] _T_2634; // @[Bitwise.scala 48:55:@1990.4]
  wire [1:0] _GEN_586; // @[Bitwise.scala 48:55:@1991.4]
  wire [2:0] _T_2635; // @[Bitwise.scala 48:55:@1991.4]
  wire [2:0] _GEN_587; // @[Bitwise.scala 48:55:@1992.4]
  wire [3:0] _T_2636; // @[Bitwise.scala 48:55:@1992.4]
  wire [4:0] _T_2637; // @[Bitwise.scala 48:55:@1993.4]
  wire [5:0] _T_2638; // @[Bitwise.scala 48:55:@1994.4]
  wire [19:0] _T_2702; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2059.4]
  wire  _T_2703; // @[Bitwise.scala 50:65:@2060.4]
  wire  _T_2704; // @[Bitwise.scala 50:65:@2061.4]
  wire  _T_2705; // @[Bitwise.scala 50:65:@2062.4]
  wire  _T_2706; // @[Bitwise.scala 50:65:@2063.4]
  wire  _T_2707; // @[Bitwise.scala 50:65:@2064.4]
  wire  _T_2708; // @[Bitwise.scala 50:65:@2065.4]
  wire  _T_2709; // @[Bitwise.scala 50:65:@2066.4]
  wire  _T_2710; // @[Bitwise.scala 50:65:@2067.4]
  wire  _T_2711; // @[Bitwise.scala 50:65:@2068.4]
  wire  _T_2712; // @[Bitwise.scala 50:65:@2069.4]
  wire  _T_2713; // @[Bitwise.scala 50:65:@2070.4]
  wire  _T_2714; // @[Bitwise.scala 50:65:@2071.4]
  wire  _T_2715; // @[Bitwise.scala 50:65:@2072.4]
  wire  _T_2716; // @[Bitwise.scala 50:65:@2073.4]
  wire  _T_2717; // @[Bitwise.scala 50:65:@2074.4]
  wire  _T_2718; // @[Bitwise.scala 50:65:@2075.4]
  wire  _T_2719; // @[Bitwise.scala 50:65:@2076.4]
  wire  _T_2720; // @[Bitwise.scala 50:65:@2077.4]
  wire  _T_2721; // @[Bitwise.scala 50:65:@2078.4]
  wire  _T_2722; // @[Bitwise.scala 50:65:@2079.4]
  wire [1:0] _T_2723; // @[Bitwise.scala 48:55:@2080.4]
  wire [1:0] _T_2724; // @[Bitwise.scala 48:55:@2081.4]
  wire [1:0] _GEN_588; // @[Bitwise.scala 48:55:@2082.4]
  wire [2:0] _T_2725; // @[Bitwise.scala 48:55:@2082.4]
  wire [2:0] _GEN_589; // @[Bitwise.scala 48:55:@2083.4]
  wire [3:0] _T_2726; // @[Bitwise.scala 48:55:@2083.4]
  wire [1:0] _T_2727; // @[Bitwise.scala 48:55:@2084.4]
  wire [1:0] _T_2728; // @[Bitwise.scala 48:55:@2085.4]
  wire [1:0] _GEN_590; // @[Bitwise.scala 48:55:@2086.4]
  wire [2:0] _T_2729; // @[Bitwise.scala 48:55:@2086.4]
  wire [2:0] _GEN_591; // @[Bitwise.scala 48:55:@2087.4]
  wire [3:0] _T_2730; // @[Bitwise.scala 48:55:@2087.4]
  wire [4:0] _T_2731; // @[Bitwise.scala 48:55:@2088.4]
  wire [1:0] _T_2732; // @[Bitwise.scala 48:55:@2089.4]
  wire [1:0] _T_2733; // @[Bitwise.scala 48:55:@2090.4]
  wire [1:0] _GEN_592; // @[Bitwise.scala 48:55:@2091.4]
  wire [2:0] _T_2734; // @[Bitwise.scala 48:55:@2091.4]
  wire [2:0] _GEN_593; // @[Bitwise.scala 48:55:@2092.4]
  wire [3:0] _T_2735; // @[Bitwise.scala 48:55:@2092.4]
  wire [1:0] _T_2736; // @[Bitwise.scala 48:55:@2093.4]
  wire [1:0] _T_2737; // @[Bitwise.scala 48:55:@2094.4]
  wire [1:0] _GEN_594; // @[Bitwise.scala 48:55:@2095.4]
  wire [2:0] _T_2738; // @[Bitwise.scala 48:55:@2095.4]
  wire [2:0] _GEN_595; // @[Bitwise.scala 48:55:@2096.4]
  wire [3:0] _T_2739; // @[Bitwise.scala 48:55:@2096.4]
  wire [4:0] _T_2740; // @[Bitwise.scala 48:55:@2097.4]
  wire [5:0] _T_2741; // @[Bitwise.scala 48:55:@2098.4]
  wire [20:0] _T_2805; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2163.4]
  wire  _T_2806; // @[Bitwise.scala 50:65:@2164.4]
  wire  _T_2807; // @[Bitwise.scala 50:65:@2165.4]
  wire  _T_2808; // @[Bitwise.scala 50:65:@2166.4]
  wire  _T_2809; // @[Bitwise.scala 50:65:@2167.4]
  wire  _T_2810; // @[Bitwise.scala 50:65:@2168.4]
  wire  _T_2811; // @[Bitwise.scala 50:65:@2169.4]
  wire  _T_2812; // @[Bitwise.scala 50:65:@2170.4]
  wire  _T_2813; // @[Bitwise.scala 50:65:@2171.4]
  wire  _T_2814; // @[Bitwise.scala 50:65:@2172.4]
  wire  _T_2815; // @[Bitwise.scala 50:65:@2173.4]
  wire  _T_2816; // @[Bitwise.scala 50:65:@2174.4]
  wire  _T_2817; // @[Bitwise.scala 50:65:@2175.4]
  wire  _T_2818; // @[Bitwise.scala 50:65:@2176.4]
  wire  _T_2819; // @[Bitwise.scala 50:65:@2177.4]
  wire  _T_2820; // @[Bitwise.scala 50:65:@2178.4]
  wire  _T_2821; // @[Bitwise.scala 50:65:@2179.4]
  wire  _T_2822; // @[Bitwise.scala 50:65:@2180.4]
  wire  _T_2823; // @[Bitwise.scala 50:65:@2181.4]
  wire  _T_2824; // @[Bitwise.scala 50:65:@2182.4]
  wire  _T_2825; // @[Bitwise.scala 50:65:@2183.4]
  wire  _T_2826; // @[Bitwise.scala 50:65:@2184.4]
  wire [1:0] _T_2827; // @[Bitwise.scala 48:55:@2185.4]
  wire [1:0] _T_2828; // @[Bitwise.scala 48:55:@2186.4]
  wire [1:0] _GEN_596; // @[Bitwise.scala 48:55:@2187.4]
  wire [2:0] _T_2829; // @[Bitwise.scala 48:55:@2187.4]
  wire [2:0] _GEN_597; // @[Bitwise.scala 48:55:@2188.4]
  wire [3:0] _T_2830; // @[Bitwise.scala 48:55:@2188.4]
  wire [1:0] _T_2831; // @[Bitwise.scala 48:55:@2189.4]
  wire [1:0] _T_2832; // @[Bitwise.scala 48:55:@2190.4]
  wire [1:0] _GEN_598; // @[Bitwise.scala 48:55:@2191.4]
  wire [2:0] _T_2833; // @[Bitwise.scala 48:55:@2191.4]
  wire [2:0] _GEN_599; // @[Bitwise.scala 48:55:@2192.4]
  wire [3:0] _T_2834; // @[Bitwise.scala 48:55:@2192.4]
  wire [4:0] _T_2835; // @[Bitwise.scala 48:55:@2193.4]
  wire [1:0] _T_2836; // @[Bitwise.scala 48:55:@2194.4]
  wire [1:0] _T_2837; // @[Bitwise.scala 48:55:@2195.4]
  wire [1:0] _GEN_600; // @[Bitwise.scala 48:55:@2196.4]
  wire [2:0] _T_2838; // @[Bitwise.scala 48:55:@2196.4]
  wire [2:0] _GEN_601; // @[Bitwise.scala 48:55:@2197.4]
  wire [3:0] _T_2839; // @[Bitwise.scala 48:55:@2197.4]
  wire [1:0] _T_2840; // @[Bitwise.scala 48:55:@2198.4]
  wire [1:0] _GEN_602; // @[Bitwise.scala 48:55:@2199.4]
  wire [2:0] _T_2841; // @[Bitwise.scala 48:55:@2199.4]
  wire [1:0] _T_2842; // @[Bitwise.scala 48:55:@2200.4]
  wire [1:0] _GEN_603; // @[Bitwise.scala 48:55:@2201.4]
  wire [2:0] _T_2843; // @[Bitwise.scala 48:55:@2201.4]
  wire [3:0] _T_2844; // @[Bitwise.scala 48:55:@2202.4]
  wire [4:0] _T_2845; // @[Bitwise.scala 48:55:@2203.4]
  wire [5:0] _T_2846; // @[Bitwise.scala 48:55:@2204.4]
  wire [21:0] _T_2910; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2269.4]
  wire  _T_2911; // @[Bitwise.scala 50:65:@2270.4]
  wire  _T_2912; // @[Bitwise.scala 50:65:@2271.4]
  wire  _T_2913; // @[Bitwise.scala 50:65:@2272.4]
  wire  _T_2914; // @[Bitwise.scala 50:65:@2273.4]
  wire  _T_2915; // @[Bitwise.scala 50:65:@2274.4]
  wire  _T_2916; // @[Bitwise.scala 50:65:@2275.4]
  wire  _T_2917; // @[Bitwise.scala 50:65:@2276.4]
  wire  _T_2918; // @[Bitwise.scala 50:65:@2277.4]
  wire  _T_2919; // @[Bitwise.scala 50:65:@2278.4]
  wire  _T_2920; // @[Bitwise.scala 50:65:@2279.4]
  wire  _T_2921; // @[Bitwise.scala 50:65:@2280.4]
  wire  _T_2922; // @[Bitwise.scala 50:65:@2281.4]
  wire  _T_2923; // @[Bitwise.scala 50:65:@2282.4]
  wire  _T_2924; // @[Bitwise.scala 50:65:@2283.4]
  wire  _T_2925; // @[Bitwise.scala 50:65:@2284.4]
  wire  _T_2926; // @[Bitwise.scala 50:65:@2285.4]
  wire  _T_2927; // @[Bitwise.scala 50:65:@2286.4]
  wire  _T_2928; // @[Bitwise.scala 50:65:@2287.4]
  wire  _T_2929; // @[Bitwise.scala 50:65:@2288.4]
  wire  _T_2930; // @[Bitwise.scala 50:65:@2289.4]
  wire  _T_2931; // @[Bitwise.scala 50:65:@2290.4]
  wire  _T_2932; // @[Bitwise.scala 50:65:@2291.4]
  wire [1:0] _T_2933; // @[Bitwise.scala 48:55:@2292.4]
  wire [1:0] _T_2934; // @[Bitwise.scala 48:55:@2293.4]
  wire [1:0] _GEN_604; // @[Bitwise.scala 48:55:@2294.4]
  wire [2:0] _T_2935; // @[Bitwise.scala 48:55:@2294.4]
  wire [2:0] _GEN_605; // @[Bitwise.scala 48:55:@2295.4]
  wire [3:0] _T_2936; // @[Bitwise.scala 48:55:@2295.4]
  wire [1:0] _T_2937; // @[Bitwise.scala 48:55:@2296.4]
  wire [1:0] _GEN_606; // @[Bitwise.scala 48:55:@2297.4]
  wire [2:0] _T_2938; // @[Bitwise.scala 48:55:@2297.4]
  wire [1:0] _T_2939; // @[Bitwise.scala 48:55:@2298.4]
  wire [1:0] _GEN_607; // @[Bitwise.scala 48:55:@2299.4]
  wire [2:0] _T_2940; // @[Bitwise.scala 48:55:@2299.4]
  wire [3:0] _T_2941; // @[Bitwise.scala 48:55:@2300.4]
  wire [4:0] _T_2942; // @[Bitwise.scala 48:55:@2301.4]
  wire [1:0] _T_2943; // @[Bitwise.scala 48:55:@2302.4]
  wire [1:0] _T_2944; // @[Bitwise.scala 48:55:@2303.4]
  wire [1:0] _GEN_608; // @[Bitwise.scala 48:55:@2304.4]
  wire [2:0] _T_2945; // @[Bitwise.scala 48:55:@2304.4]
  wire [2:0] _GEN_609; // @[Bitwise.scala 48:55:@2305.4]
  wire [3:0] _T_2946; // @[Bitwise.scala 48:55:@2305.4]
  wire [1:0] _T_2947; // @[Bitwise.scala 48:55:@2306.4]
  wire [1:0] _GEN_610; // @[Bitwise.scala 48:55:@2307.4]
  wire [2:0] _T_2948; // @[Bitwise.scala 48:55:@2307.4]
  wire [1:0] _T_2949; // @[Bitwise.scala 48:55:@2308.4]
  wire [1:0] _GEN_611; // @[Bitwise.scala 48:55:@2309.4]
  wire [2:0] _T_2950; // @[Bitwise.scala 48:55:@2309.4]
  wire [3:0] _T_2951; // @[Bitwise.scala 48:55:@2310.4]
  wire [4:0] _T_2952; // @[Bitwise.scala 48:55:@2311.4]
  wire [5:0] _T_2953; // @[Bitwise.scala 48:55:@2312.4]
  wire [22:0] _T_3017; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2377.4]
  wire  _T_3018; // @[Bitwise.scala 50:65:@2378.4]
  wire  _T_3019; // @[Bitwise.scala 50:65:@2379.4]
  wire  _T_3020; // @[Bitwise.scala 50:65:@2380.4]
  wire  _T_3021; // @[Bitwise.scala 50:65:@2381.4]
  wire  _T_3022; // @[Bitwise.scala 50:65:@2382.4]
  wire  _T_3023; // @[Bitwise.scala 50:65:@2383.4]
  wire  _T_3024; // @[Bitwise.scala 50:65:@2384.4]
  wire  _T_3025; // @[Bitwise.scala 50:65:@2385.4]
  wire  _T_3026; // @[Bitwise.scala 50:65:@2386.4]
  wire  _T_3027; // @[Bitwise.scala 50:65:@2387.4]
  wire  _T_3028; // @[Bitwise.scala 50:65:@2388.4]
  wire  _T_3029; // @[Bitwise.scala 50:65:@2389.4]
  wire  _T_3030; // @[Bitwise.scala 50:65:@2390.4]
  wire  _T_3031; // @[Bitwise.scala 50:65:@2391.4]
  wire  _T_3032; // @[Bitwise.scala 50:65:@2392.4]
  wire  _T_3033; // @[Bitwise.scala 50:65:@2393.4]
  wire  _T_3034; // @[Bitwise.scala 50:65:@2394.4]
  wire  _T_3035; // @[Bitwise.scala 50:65:@2395.4]
  wire  _T_3036; // @[Bitwise.scala 50:65:@2396.4]
  wire  _T_3037; // @[Bitwise.scala 50:65:@2397.4]
  wire  _T_3038; // @[Bitwise.scala 50:65:@2398.4]
  wire  _T_3039; // @[Bitwise.scala 50:65:@2399.4]
  wire  _T_3040; // @[Bitwise.scala 50:65:@2400.4]
  wire [1:0] _T_3041; // @[Bitwise.scala 48:55:@2401.4]
  wire [1:0] _T_3042; // @[Bitwise.scala 48:55:@2402.4]
  wire [1:0] _GEN_612; // @[Bitwise.scala 48:55:@2403.4]
  wire [2:0] _T_3043; // @[Bitwise.scala 48:55:@2403.4]
  wire [2:0] _GEN_613; // @[Bitwise.scala 48:55:@2404.4]
  wire [3:0] _T_3044; // @[Bitwise.scala 48:55:@2404.4]
  wire [1:0] _T_3045; // @[Bitwise.scala 48:55:@2405.4]
  wire [1:0] _GEN_614; // @[Bitwise.scala 48:55:@2406.4]
  wire [2:0] _T_3046; // @[Bitwise.scala 48:55:@2406.4]
  wire [1:0] _T_3047; // @[Bitwise.scala 48:55:@2407.4]
  wire [1:0] _GEN_615; // @[Bitwise.scala 48:55:@2408.4]
  wire [2:0] _T_3048; // @[Bitwise.scala 48:55:@2408.4]
  wire [3:0] _T_3049; // @[Bitwise.scala 48:55:@2409.4]
  wire [4:0] _T_3050; // @[Bitwise.scala 48:55:@2410.4]
  wire [1:0] _T_3051; // @[Bitwise.scala 48:55:@2411.4]
  wire [1:0] _GEN_616; // @[Bitwise.scala 48:55:@2412.4]
  wire [2:0] _T_3052; // @[Bitwise.scala 48:55:@2412.4]
  wire [1:0] _T_3053; // @[Bitwise.scala 48:55:@2413.4]
  wire [1:0] _GEN_617; // @[Bitwise.scala 48:55:@2414.4]
  wire [2:0] _T_3054; // @[Bitwise.scala 48:55:@2414.4]
  wire [3:0] _T_3055; // @[Bitwise.scala 48:55:@2415.4]
  wire [1:0] _T_3056; // @[Bitwise.scala 48:55:@2416.4]
  wire [1:0] _GEN_618; // @[Bitwise.scala 48:55:@2417.4]
  wire [2:0] _T_3057; // @[Bitwise.scala 48:55:@2417.4]
  wire [1:0] _T_3058; // @[Bitwise.scala 48:55:@2418.4]
  wire [1:0] _GEN_619; // @[Bitwise.scala 48:55:@2419.4]
  wire [2:0] _T_3059; // @[Bitwise.scala 48:55:@2419.4]
  wire [3:0] _T_3060; // @[Bitwise.scala 48:55:@2420.4]
  wire [4:0] _T_3061; // @[Bitwise.scala 48:55:@2421.4]
  wire [5:0] _T_3062; // @[Bitwise.scala 48:55:@2422.4]
  wire [23:0] _T_3126; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2487.4]
  wire  _T_3127; // @[Bitwise.scala 50:65:@2488.4]
  wire  _T_3128; // @[Bitwise.scala 50:65:@2489.4]
  wire  _T_3129; // @[Bitwise.scala 50:65:@2490.4]
  wire  _T_3130; // @[Bitwise.scala 50:65:@2491.4]
  wire  _T_3131; // @[Bitwise.scala 50:65:@2492.4]
  wire  _T_3132; // @[Bitwise.scala 50:65:@2493.4]
  wire  _T_3133; // @[Bitwise.scala 50:65:@2494.4]
  wire  _T_3134; // @[Bitwise.scala 50:65:@2495.4]
  wire  _T_3135; // @[Bitwise.scala 50:65:@2496.4]
  wire  _T_3136; // @[Bitwise.scala 50:65:@2497.4]
  wire  _T_3137; // @[Bitwise.scala 50:65:@2498.4]
  wire  _T_3138; // @[Bitwise.scala 50:65:@2499.4]
  wire  _T_3139; // @[Bitwise.scala 50:65:@2500.4]
  wire  _T_3140; // @[Bitwise.scala 50:65:@2501.4]
  wire  _T_3141; // @[Bitwise.scala 50:65:@2502.4]
  wire  _T_3142; // @[Bitwise.scala 50:65:@2503.4]
  wire  _T_3143; // @[Bitwise.scala 50:65:@2504.4]
  wire  _T_3144; // @[Bitwise.scala 50:65:@2505.4]
  wire  _T_3145; // @[Bitwise.scala 50:65:@2506.4]
  wire  _T_3146; // @[Bitwise.scala 50:65:@2507.4]
  wire  _T_3147; // @[Bitwise.scala 50:65:@2508.4]
  wire  _T_3148; // @[Bitwise.scala 50:65:@2509.4]
  wire  _T_3149; // @[Bitwise.scala 50:65:@2510.4]
  wire  _T_3150; // @[Bitwise.scala 50:65:@2511.4]
  wire [1:0] _T_3151; // @[Bitwise.scala 48:55:@2512.4]
  wire [1:0] _GEN_620; // @[Bitwise.scala 48:55:@2513.4]
  wire [2:0] _T_3152; // @[Bitwise.scala 48:55:@2513.4]
  wire [1:0] _T_3153; // @[Bitwise.scala 48:55:@2514.4]
  wire [1:0] _GEN_621; // @[Bitwise.scala 48:55:@2515.4]
  wire [2:0] _T_3154; // @[Bitwise.scala 48:55:@2515.4]
  wire [3:0] _T_3155; // @[Bitwise.scala 48:55:@2516.4]
  wire [1:0] _T_3156; // @[Bitwise.scala 48:55:@2517.4]
  wire [1:0] _GEN_622; // @[Bitwise.scala 48:55:@2518.4]
  wire [2:0] _T_3157; // @[Bitwise.scala 48:55:@2518.4]
  wire [1:0] _T_3158; // @[Bitwise.scala 48:55:@2519.4]
  wire [1:0] _GEN_623; // @[Bitwise.scala 48:55:@2520.4]
  wire [2:0] _T_3159; // @[Bitwise.scala 48:55:@2520.4]
  wire [3:0] _T_3160; // @[Bitwise.scala 48:55:@2521.4]
  wire [4:0] _T_3161; // @[Bitwise.scala 48:55:@2522.4]
  wire [1:0] _T_3162; // @[Bitwise.scala 48:55:@2523.4]
  wire [1:0] _GEN_624; // @[Bitwise.scala 48:55:@2524.4]
  wire [2:0] _T_3163; // @[Bitwise.scala 48:55:@2524.4]
  wire [1:0] _T_3164; // @[Bitwise.scala 48:55:@2525.4]
  wire [1:0] _GEN_625; // @[Bitwise.scala 48:55:@2526.4]
  wire [2:0] _T_3165; // @[Bitwise.scala 48:55:@2526.4]
  wire [3:0] _T_3166; // @[Bitwise.scala 48:55:@2527.4]
  wire [1:0] _T_3167; // @[Bitwise.scala 48:55:@2528.4]
  wire [1:0] _GEN_626; // @[Bitwise.scala 48:55:@2529.4]
  wire [2:0] _T_3168; // @[Bitwise.scala 48:55:@2529.4]
  wire [1:0] _T_3169; // @[Bitwise.scala 48:55:@2530.4]
  wire [1:0] _GEN_627; // @[Bitwise.scala 48:55:@2531.4]
  wire [2:0] _T_3170; // @[Bitwise.scala 48:55:@2531.4]
  wire [3:0] _T_3171; // @[Bitwise.scala 48:55:@2532.4]
  wire [4:0] _T_3172; // @[Bitwise.scala 48:55:@2533.4]
  wire [5:0] _T_3173; // @[Bitwise.scala 48:55:@2534.4]
  wire [24:0] _T_3237; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2599.4]
  wire  _T_3238; // @[Bitwise.scala 50:65:@2600.4]
  wire  _T_3239; // @[Bitwise.scala 50:65:@2601.4]
  wire  _T_3240; // @[Bitwise.scala 50:65:@2602.4]
  wire  _T_3241; // @[Bitwise.scala 50:65:@2603.4]
  wire  _T_3242; // @[Bitwise.scala 50:65:@2604.4]
  wire  _T_3243; // @[Bitwise.scala 50:65:@2605.4]
  wire  _T_3244; // @[Bitwise.scala 50:65:@2606.4]
  wire  _T_3245; // @[Bitwise.scala 50:65:@2607.4]
  wire  _T_3246; // @[Bitwise.scala 50:65:@2608.4]
  wire  _T_3247; // @[Bitwise.scala 50:65:@2609.4]
  wire  _T_3248; // @[Bitwise.scala 50:65:@2610.4]
  wire  _T_3249; // @[Bitwise.scala 50:65:@2611.4]
  wire  _T_3250; // @[Bitwise.scala 50:65:@2612.4]
  wire  _T_3251; // @[Bitwise.scala 50:65:@2613.4]
  wire  _T_3252; // @[Bitwise.scala 50:65:@2614.4]
  wire  _T_3253; // @[Bitwise.scala 50:65:@2615.4]
  wire  _T_3254; // @[Bitwise.scala 50:65:@2616.4]
  wire  _T_3255; // @[Bitwise.scala 50:65:@2617.4]
  wire  _T_3256; // @[Bitwise.scala 50:65:@2618.4]
  wire  _T_3257; // @[Bitwise.scala 50:65:@2619.4]
  wire  _T_3258; // @[Bitwise.scala 50:65:@2620.4]
  wire  _T_3259; // @[Bitwise.scala 50:65:@2621.4]
  wire  _T_3260; // @[Bitwise.scala 50:65:@2622.4]
  wire  _T_3261; // @[Bitwise.scala 50:65:@2623.4]
  wire  _T_3262; // @[Bitwise.scala 50:65:@2624.4]
  wire [1:0] _T_3263; // @[Bitwise.scala 48:55:@2625.4]
  wire [1:0] _GEN_628; // @[Bitwise.scala 48:55:@2626.4]
  wire [2:0] _T_3264; // @[Bitwise.scala 48:55:@2626.4]
  wire [1:0] _T_3265; // @[Bitwise.scala 48:55:@2627.4]
  wire [1:0] _GEN_629; // @[Bitwise.scala 48:55:@2628.4]
  wire [2:0] _T_3266; // @[Bitwise.scala 48:55:@2628.4]
  wire [3:0] _T_3267; // @[Bitwise.scala 48:55:@2629.4]
  wire [1:0] _T_3268; // @[Bitwise.scala 48:55:@2630.4]
  wire [1:0] _GEN_630; // @[Bitwise.scala 48:55:@2631.4]
  wire [2:0] _T_3269; // @[Bitwise.scala 48:55:@2631.4]
  wire [1:0] _T_3270; // @[Bitwise.scala 48:55:@2632.4]
  wire [1:0] _GEN_631; // @[Bitwise.scala 48:55:@2633.4]
  wire [2:0] _T_3271; // @[Bitwise.scala 48:55:@2633.4]
  wire [3:0] _T_3272; // @[Bitwise.scala 48:55:@2634.4]
  wire [4:0] _T_3273; // @[Bitwise.scala 48:55:@2635.4]
  wire [1:0] _T_3274; // @[Bitwise.scala 48:55:@2636.4]
  wire [1:0] _GEN_632; // @[Bitwise.scala 48:55:@2637.4]
  wire [2:0] _T_3275; // @[Bitwise.scala 48:55:@2637.4]
  wire [1:0] _T_3276; // @[Bitwise.scala 48:55:@2638.4]
  wire [1:0] _GEN_633; // @[Bitwise.scala 48:55:@2639.4]
  wire [2:0] _T_3277; // @[Bitwise.scala 48:55:@2639.4]
  wire [3:0] _T_3278; // @[Bitwise.scala 48:55:@2640.4]
  wire [1:0] _T_3279; // @[Bitwise.scala 48:55:@2641.4]
  wire [1:0] _GEN_634; // @[Bitwise.scala 48:55:@2642.4]
  wire [2:0] _T_3280; // @[Bitwise.scala 48:55:@2642.4]
  wire [1:0] _T_3281; // @[Bitwise.scala 48:55:@2643.4]
  wire [1:0] _T_3282; // @[Bitwise.scala 48:55:@2644.4]
  wire [2:0] _T_3283; // @[Bitwise.scala 48:55:@2645.4]
  wire [3:0] _T_3284; // @[Bitwise.scala 48:55:@2646.4]
  wire [4:0] _T_3285; // @[Bitwise.scala 48:55:@2647.4]
  wire [5:0] _T_3286; // @[Bitwise.scala 48:55:@2648.4]
  wire [25:0] _T_3350; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2713.4]
  wire  _T_3351; // @[Bitwise.scala 50:65:@2714.4]
  wire  _T_3352; // @[Bitwise.scala 50:65:@2715.4]
  wire  _T_3353; // @[Bitwise.scala 50:65:@2716.4]
  wire  _T_3354; // @[Bitwise.scala 50:65:@2717.4]
  wire  _T_3355; // @[Bitwise.scala 50:65:@2718.4]
  wire  _T_3356; // @[Bitwise.scala 50:65:@2719.4]
  wire  _T_3357; // @[Bitwise.scala 50:65:@2720.4]
  wire  _T_3358; // @[Bitwise.scala 50:65:@2721.4]
  wire  _T_3359; // @[Bitwise.scala 50:65:@2722.4]
  wire  _T_3360; // @[Bitwise.scala 50:65:@2723.4]
  wire  _T_3361; // @[Bitwise.scala 50:65:@2724.4]
  wire  _T_3362; // @[Bitwise.scala 50:65:@2725.4]
  wire  _T_3363; // @[Bitwise.scala 50:65:@2726.4]
  wire  _T_3364; // @[Bitwise.scala 50:65:@2727.4]
  wire  _T_3365; // @[Bitwise.scala 50:65:@2728.4]
  wire  _T_3366; // @[Bitwise.scala 50:65:@2729.4]
  wire  _T_3367; // @[Bitwise.scala 50:65:@2730.4]
  wire  _T_3368; // @[Bitwise.scala 50:65:@2731.4]
  wire  _T_3369; // @[Bitwise.scala 50:65:@2732.4]
  wire  _T_3370; // @[Bitwise.scala 50:65:@2733.4]
  wire  _T_3371; // @[Bitwise.scala 50:65:@2734.4]
  wire  _T_3372; // @[Bitwise.scala 50:65:@2735.4]
  wire  _T_3373; // @[Bitwise.scala 50:65:@2736.4]
  wire  _T_3374; // @[Bitwise.scala 50:65:@2737.4]
  wire  _T_3375; // @[Bitwise.scala 50:65:@2738.4]
  wire  _T_3376; // @[Bitwise.scala 50:65:@2739.4]
  wire [1:0] _T_3377; // @[Bitwise.scala 48:55:@2740.4]
  wire [1:0] _GEN_635; // @[Bitwise.scala 48:55:@2741.4]
  wire [2:0] _T_3378; // @[Bitwise.scala 48:55:@2741.4]
  wire [1:0] _T_3379; // @[Bitwise.scala 48:55:@2742.4]
  wire [1:0] _GEN_636; // @[Bitwise.scala 48:55:@2743.4]
  wire [2:0] _T_3380; // @[Bitwise.scala 48:55:@2743.4]
  wire [3:0] _T_3381; // @[Bitwise.scala 48:55:@2744.4]
  wire [1:0] _T_3382; // @[Bitwise.scala 48:55:@2745.4]
  wire [1:0] _GEN_637; // @[Bitwise.scala 48:55:@2746.4]
  wire [2:0] _T_3383; // @[Bitwise.scala 48:55:@2746.4]
  wire [1:0] _T_3384; // @[Bitwise.scala 48:55:@2747.4]
  wire [1:0] _T_3385; // @[Bitwise.scala 48:55:@2748.4]
  wire [2:0] _T_3386; // @[Bitwise.scala 48:55:@2749.4]
  wire [3:0] _T_3387; // @[Bitwise.scala 48:55:@2750.4]
  wire [4:0] _T_3388; // @[Bitwise.scala 48:55:@2751.4]
  wire [1:0] _T_3389; // @[Bitwise.scala 48:55:@2752.4]
  wire [1:0] _GEN_638; // @[Bitwise.scala 48:55:@2753.4]
  wire [2:0] _T_3390; // @[Bitwise.scala 48:55:@2753.4]
  wire [1:0] _T_3391; // @[Bitwise.scala 48:55:@2754.4]
  wire [1:0] _GEN_639; // @[Bitwise.scala 48:55:@2755.4]
  wire [2:0] _T_3392; // @[Bitwise.scala 48:55:@2755.4]
  wire [3:0] _T_3393; // @[Bitwise.scala 48:55:@2756.4]
  wire [1:0] _T_3394; // @[Bitwise.scala 48:55:@2757.4]
  wire [1:0] _GEN_640; // @[Bitwise.scala 48:55:@2758.4]
  wire [2:0] _T_3395; // @[Bitwise.scala 48:55:@2758.4]
  wire [1:0] _T_3396; // @[Bitwise.scala 48:55:@2759.4]
  wire [1:0] _T_3397; // @[Bitwise.scala 48:55:@2760.4]
  wire [2:0] _T_3398; // @[Bitwise.scala 48:55:@2761.4]
  wire [3:0] _T_3399; // @[Bitwise.scala 48:55:@2762.4]
  wire [4:0] _T_3400; // @[Bitwise.scala 48:55:@2763.4]
  wire [5:0] _T_3401; // @[Bitwise.scala 48:55:@2764.4]
  wire [26:0] _T_3465; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2829.4]
  wire  _T_3466; // @[Bitwise.scala 50:65:@2830.4]
  wire  _T_3467; // @[Bitwise.scala 50:65:@2831.4]
  wire  _T_3468; // @[Bitwise.scala 50:65:@2832.4]
  wire  _T_3469; // @[Bitwise.scala 50:65:@2833.4]
  wire  _T_3470; // @[Bitwise.scala 50:65:@2834.4]
  wire  _T_3471; // @[Bitwise.scala 50:65:@2835.4]
  wire  _T_3472; // @[Bitwise.scala 50:65:@2836.4]
  wire  _T_3473; // @[Bitwise.scala 50:65:@2837.4]
  wire  _T_3474; // @[Bitwise.scala 50:65:@2838.4]
  wire  _T_3475; // @[Bitwise.scala 50:65:@2839.4]
  wire  _T_3476; // @[Bitwise.scala 50:65:@2840.4]
  wire  _T_3477; // @[Bitwise.scala 50:65:@2841.4]
  wire  _T_3478; // @[Bitwise.scala 50:65:@2842.4]
  wire  _T_3479; // @[Bitwise.scala 50:65:@2843.4]
  wire  _T_3480; // @[Bitwise.scala 50:65:@2844.4]
  wire  _T_3481; // @[Bitwise.scala 50:65:@2845.4]
  wire  _T_3482; // @[Bitwise.scala 50:65:@2846.4]
  wire  _T_3483; // @[Bitwise.scala 50:65:@2847.4]
  wire  _T_3484; // @[Bitwise.scala 50:65:@2848.4]
  wire  _T_3485; // @[Bitwise.scala 50:65:@2849.4]
  wire  _T_3486; // @[Bitwise.scala 50:65:@2850.4]
  wire  _T_3487; // @[Bitwise.scala 50:65:@2851.4]
  wire  _T_3488; // @[Bitwise.scala 50:65:@2852.4]
  wire  _T_3489; // @[Bitwise.scala 50:65:@2853.4]
  wire  _T_3490; // @[Bitwise.scala 50:65:@2854.4]
  wire  _T_3491; // @[Bitwise.scala 50:65:@2855.4]
  wire  _T_3492; // @[Bitwise.scala 50:65:@2856.4]
  wire [1:0] _T_3493; // @[Bitwise.scala 48:55:@2857.4]
  wire [1:0] _GEN_641; // @[Bitwise.scala 48:55:@2858.4]
  wire [2:0] _T_3494; // @[Bitwise.scala 48:55:@2858.4]
  wire [1:0] _T_3495; // @[Bitwise.scala 48:55:@2859.4]
  wire [1:0] _GEN_642; // @[Bitwise.scala 48:55:@2860.4]
  wire [2:0] _T_3496; // @[Bitwise.scala 48:55:@2860.4]
  wire [3:0] _T_3497; // @[Bitwise.scala 48:55:@2861.4]
  wire [1:0] _T_3498; // @[Bitwise.scala 48:55:@2862.4]
  wire [1:0] _GEN_643; // @[Bitwise.scala 48:55:@2863.4]
  wire [2:0] _T_3499; // @[Bitwise.scala 48:55:@2863.4]
  wire [1:0] _T_3500; // @[Bitwise.scala 48:55:@2864.4]
  wire [1:0] _T_3501; // @[Bitwise.scala 48:55:@2865.4]
  wire [2:0] _T_3502; // @[Bitwise.scala 48:55:@2866.4]
  wire [3:0] _T_3503; // @[Bitwise.scala 48:55:@2867.4]
  wire [4:0] _T_3504; // @[Bitwise.scala 48:55:@2868.4]
  wire [1:0] _T_3505; // @[Bitwise.scala 48:55:@2869.4]
  wire [1:0] _GEN_644; // @[Bitwise.scala 48:55:@2870.4]
  wire [2:0] _T_3506; // @[Bitwise.scala 48:55:@2870.4]
  wire [1:0] _T_3507; // @[Bitwise.scala 48:55:@2871.4]
  wire [1:0] _T_3508; // @[Bitwise.scala 48:55:@2872.4]
  wire [2:0] _T_3509; // @[Bitwise.scala 48:55:@2873.4]
  wire [3:0] _T_3510; // @[Bitwise.scala 48:55:@2874.4]
  wire [1:0] _T_3511; // @[Bitwise.scala 48:55:@2875.4]
  wire [1:0] _GEN_645; // @[Bitwise.scala 48:55:@2876.4]
  wire [2:0] _T_3512; // @[Bitwise.scala 48:55:@2876.4]
  wire [1:0] _T_3513; // @[Bitwise.scala 48:55:@2877.4]
  wire [1:0] _T_3514; // @[Bitwise.scala 48:55:@2878.4]
  wire [2:0] _T_3515; // @[Bitwise.scala 48:55:@2879.4]
  wire [3:0] _T_3516; // @[Bitwise.scala 48:55:@2880.4]
  wire [4:0] _T_3517; // @[Bitwise.scala 48:55:@2881.4]
  wire [5:0] _T_3518; // @[Bitwise.scala 48:55:@2882.4]
  wire [27:0] _T_3582; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2947.4]
  wire  _T_3583; // @[Bitwise.scala 50:65:@2948.4]
  wire  _T_3584; // @[Bitwise.scala 50:65:@2949.4]
  wire  _T_3585; // @[Bitwise.scala 50:65:@2950.4]
  wire  _T_3586; // @[Bitwise.scala 50:65:@2951.4]
  wire  _T_3587; // @[Bitwise.scala 50:65:@2952.4]
  wire  _T_3588; // @[Bitwise.scala 50:65:@2953.4]
  wire  _T_3589; // @[Bitwise.scala 50:65:@2954.4]
  wire  _T_3590; // @[Bitwise.scala 50:65:@2955.4]
  wire  _T_3591; // @[Bitwise.scala 50:65:@2956.4]
  wire  _T_3592; // @[Bitwise.scala 50:65:@2957.4]
  wire  _T_3593; // @[Bitwise.scala 50:65:@2958.4]
  wire  _T_3594; // @[Bitwise.scala 50:65:@2959.4]
  wire  _T_3595; // @[Bitwise.scala 50:65:@2960.4]
  wire  _T_3596; // @[Bitwise.scala 50:65:@2961.4]
  wire  _T_3597; // @[Bitwise.scala 50:65:@2962.4]
  wire  _T_3598; // @[Bitwise.scala 50:65:@2963.4]
  wire  _T_3599; // @[Bitwise.scala 50:65:@2964.4]
  wire  _T_3600; // @[Bitwise.scala 50:65:@2965.4]
  wire  _T_3601; // @[Bitwise.scala 50:65:@2966.4]
  wire  _T_3602; // @[Bitwise.scala 50:65:@2967.4]
  wire  _T_3603; // @[Bitwise.scala 50:65:@2968.4]
  wire  _T_3604; // @[Bitwise.scala 50:65:@2969.4]
  wire  _T_3605; // @[Bitwise.scala 50:65:@2970.4]
  wire  _T_3606; // @[Bitwise.scala 50:65:@2971.4]
  wire  _T_3607; // @[Bitwise.scala 50:65:@2972.4]
  wire  _T_3608; // @[Bitwise.scala 50:65:@2973.4]
  wire  _T_3609; // @[Bitwise.scala 50:65:@2974.4]
  wire  _T_3610; // @[Bitwise.scala 50:65:@2975.4]
  wire [1:0] _T_3611; // @[Bitwise.scala 48:55:@2976.4]
  wire [1:0] _GEN_646; // @[Bitwise.scala 48:55:@2977.4]
  wire [2:0] _T_3612; // @[Bitwise.scala 48:55:@2977.4]
  wire [1:0] _T_3613; // @[Bitwise.scala 48:55:@2978.4]
  wire [1:0] _T_3614; // @[Bitwise.scala 48:55:@2979.4]
  wire [2:0] _T_3615; // @[Bitwise.scala 48:55:@2980.4]
  wire [3:0] _T_3616; // @[Bitwise.scala 48:55:@2981.4]
  wire [1:0] _T_3617; // @[Bitwise.scala 48:55:@2982.4]
  wire [1:0] _GEN_647; // @[Bitwise.scala 48:55:@2983.4]
  wire [2:0] _T_3618; // @[Bitwise.scala 48:55:@2983.4]
  wire [1:0] _T_3619; // @[Bitwise.scala 48:55:@2984.4]
  wire [1:0] _T_3620; // @[Bitwise.scala 48:55:@2985.4]
  wire [2:0] _T_3621; // @[Bitwise.scala 48:55:@2986.4]
  wire [3:0] _T_3622; // @[Bitwise.scala 48:55:@2987.4]
  wire [4:0] _T_3623; // @[Bitwise.scala 48:55:@2988.4]
  wire [1:0] _T_3624; // @[Bitwise.scala 48:55:@2989.4]
  wire [1:0] _GEN_648; // @[Bitwise.scala 48:55:@2990.4]
  wire [2:0] _T_3625; // @[Bitwise.scala 48:55:@2990.4]
  wire [1:0] _T_3626; // @[Bitwise.scala 48:55:@2991.4]
  wire [1:0] _T_3627; // @[Bitwise.scala 48:55:@2992.4]
  wire [2:0] _T_3628; // @[Bitwise.scala 48:55:@2993.4]
  wire [3:0] _T_3629; // @[Bitwise.scala 48:55:@2994.4]
  wire [1:0] _T_3630; // @[Bitwise.scala 48:55:@2995.4]
  wire [1:0] _GEN_649; // @[Bitwise.scala 48:55:@2996.4]
  wire [2:0] _T_3631; // @[Bitwise.scala 48:55:@2996.4]
  wire [1:0] _T_3632; // @[Bitwise.scala 48:55:@2997.4]
  wire [1:0] _T_3633; // @[Bitwise.scala 48:55:@2998.4]
  wire [2:0] _T_3634; // @[Bitwise.scala 48:55:@2999.4]
  wire [3:0] _T_3635; // @[Bitwise.scala 48:55:@3000.4]
  wire [4:0] _T_3636; // @[Bitwise.scala 48:55:@3001.4]
  wire [5:0] _T_3637; // @[Bitwise.scala 48:55:@3002.4]
  wire [28:0] _T_3701; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3067.4]
  wire  _T_3702; // @[Bitwise.scala 50:65:@3068.4]
  wire  _T_3703; // @[Bitwise.scala 50:65:@3069.4]
  wire  _T_3704; // @[Bitwise.scala 50:65:@3070.4]
  wire  _T_3705; // @[Bitwise.scala 50:65:@3071.4]
  wire  _T_3706; // @[Bitwise.scala 50:65:@3072.4]
  wire  _T_3707; // @[Bitwise.scala 50:65:@3073.4]
  wire  _T_3708; // @[Bitwise.scala 50:65:@3074.4]
  wire  _T_3709; // @[Bitwise.scala 50:65:@3075.4]
  wire  _T_3710; // @[Bitwise.scala 50:65:@3076.4]
  wire  _T_3711; // @[Bitwise.scala 50:65:@3077.4]
  wire  _T_3712; // @[Bitwise.scala 50:65:@3078.4]
  wire  _T_3713; // @[Bitwise.scala 50:65:@3079.4]
  wire  _T_3714; // @[Bitwise.scala 50:65:@3080.4]
  wire  _T_3715; // @[Bitwise.scala 50:65:@3081.4]
  wire  _T_3716; // @[Bitwise.scala 50:65:@3082.4]
  wire  _T_3717; // @[Bitwise.scala 50:65:@3083.4]
  wire  _T_3718; // @[Bitwise.scala 50:65:@3084.4]
  wire  _T_3719; // @[Bitwise.scala 50:65:@3085.4]
  wire  _T_3720; // @[Bitwise.scala 50:65:@3086.4]
  wire  _T_3721; // @[Bitwise.scala 50:65:@3087.4]
  wire  _T_3722; // @[Bitwise.scala 50:65:@3088.4]
  wire  _T_3723; // @[Bitwise.scala 50:65:@3089.4]
  wire  _T_3724; // @[Bitwise.scala 50:65:@3090.4]
  wire  _T_3725; // @[Bitwise.scala 50:65:@3091.4]
  wire  _T_3726; // @[Bitwise.scala 50:65:@3092.4]
  wire  _T_3727; // @[Bitwise.scala 50:65:@3093.4]
  wire  _T_3728; // @[Bitwise.scala 50:65:@3094.4]
  wire  _T_3729; // @[Bitwise.scala 50:65:@3095.4]
  wire  _T_3730; // @[Bitwise.scala 50:65:@3096.4]
  wire [1:0] _T_3731; // @[Bitwise.scala 48:55:@3097.4]
  wire [1:0] _GEN_650; // @[Bitwise.scala 48:55:@3098.4]
  wire [2:0] _T_3732; // @[Bitwise.scala 48:55:@3098.4]
  wire [1:0] _T_3733; // @[Bitwise.scala 48:55:@3099.4]
  wire [1:0] _T_3734; // @[Bitwise.scala 48:55:@3100.4]
  wire [2:0] _T_3735; // @[Bitwise.scala 48:55:@3101.4]
  wire [3:0] _T_3736; // @[Bitwise.scala 48:55:@3102.4]
  wire [1:0] _T_3737; // @[Bitwise.scala 48:55:@3103.4]
  wire [1:0] _GEN_651; // @[Bitwise.scala 48:55:@3104.4]
  wire [2:0] _T_3738; // @[Bitwise.scala 48:55:@3104.4]
  wire [1:0] _T_3739; // @[Bitwise.scala 48:55:@3105.4]
  wire [1:0] _T_3740; // @[Bitwise.scala 48:55:@3106.4]
  wire [2:0] _T_3741; // @[Bitwise.scala 48:55:@3107.4]
  wire [3:0] _T_3742; // @[Bitwise.scala 48:55:@3108.4]
  wire [4:0] _T_3743; // @[Bitwise.scala 48:55:@3109.4]
  wire [1:0] _T_3744; // @[Bitwise.scala 48:55:@3110.4]
  wire [1:0] _GEN_652; // @[Bitwise.scala 48:55:@3111.4]
  wire [2:0] _T_3745; // @[Bitwise.scala 48:55:@3111.4]
  wire [1:0] _T_3746; // @[Bitwise.scala 48:55:@3112.4]
  wire [1:0] _T_3747; // @[Bitwise.scala 48:55:@3113.4]
  wire [2:0] _T_3748; // @[Bitwise.scala 48:55:@3114.4]
  wire [3:0] _T_3749; // @[Bitwise.scala 48:55:@3115.4]
  wire [1:0] _T_3750; // @[Bitwise.scala 48:55:@3116.4]
  wire [1:0] _T_3751; // @[Bitwise.scala 48:55:@3117.4]
  wire [2:0] _T_3752; // @[Bitwise.scala 48:55:@3118.4]
  wire [1:0] _T_3753; // @[Bitwise.scala 48:55:@3119.4]
  wire [1:0] _T_3754; // @[Bitwise.scala 48:55:@3120.4]
  wire [2:0] _T_3755; // @[Bitwise.scala 48:55:@3121.4]
  wire [3:0] _T_3756; // @[Bitwise.scala 48:55:@3122.4]
  wire [4:0] _T_3757; // @[Bitwise.scala 48:55:@3123.4]
  wire [5:0] _T_3758; // @[Bitwise.scala 48:55:@3124.4]
  wire [29:0] _T_3822; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3189.4]
  wire  _T_3823; // @[Bitwise.scala 50:65:@3190.4]
  wire  _T_3824; // @[Bitwise.scala 50:65:@3191.4]
  wire  _T_3825; // @[Bitwise.scala 50:65:@3192.4]
  wire  _T_3826; // @[Bitwise.scala 50:65:@3193.4]
  wire  _T_3827; // @[Bitwise.scala 50:65:@3194.4]
  wire  _T_3828; // @[Bitwise.scala 50:65:@3195.4]
  wire  _T_3829; // @[Bitwise.scala 50:65:@3196.4]
  wire  _T_3830; // @[Bitwise.scala 50:65:@3197.4]
  wire  _T_3831; // @[Bitwise.scala 50:65:@3198.4]
  wire  _T_3832; // @[Bitwise.scala 50:65:@3199.4]
  wire  _T_3833; // @[Bitwise.scala 50:65:@3200.4]
  wire  _T_3834; // @[Bitwise.scala 50:65:@3201.4]
  wire  _T_3835; // @[Bitwise.scala 50:65:@3202.4]
  wire  _T_3836; // @[Bitwise.scala 50:65:@3203.4]
  wire  _T_3837; // @[Bitwise.scala 50:65:@3204.4]
  wire  _T_3838; // @[Bitwise.scala 50:65:@3205.4]
  wire  _T_3839; // @[Bitwise.scala 50:65:@3206.4]
  wire  _T_3840; // @[Bitwise.scala 50:65:@3207.4]
  wire  _T_3841; // @[Bitwise.scala 50:65:@3208.4]
  wire  _T_3842; // @[Bitwise.scala 50:65:@3209.4]
  wire  _T_3843; // @[Bitwise.scala 50:65:@3210.4]
  wire  _T_3844; // @[Bitwise.scala 50:65:@3211.4]
  wire  _T_3845; // @[Bitwise.scala 50:65:@3212.4]
  wire  _T_3846; // @[Bitwise.scala 50:65:@3213.4]
  wire  _T_3847; // @[Bitwise.scala 50:65:@3214.4]
  wire  _T_3848; // @[Bitwise.scala 50:65:@3215.4]
  wire  _T_3849; // @[Bitwise.scala 50:65:@3216.4]
  wire  _T_3850; // @[Bitwise.scala 50:65:@3217.4]
  wire  _T_3851; // @[Bitwise.scala 50:65:@3218.4]
  wire  _T_3852; // @[Bitwise.scala 50:65:@3219.4]
  wire [1:0] _T_3853; // @[Bitwise.scala 48:55:@3220.4]
  wire [1:0] _GEN_653; // @[Bitwise.scala 48:55:@3221.4]
  wire [2:0] _T_3854; // @[Bitwise.scala 48:55:@3221.4]
  wire [1:0] _T_3855; // @[Bitwise.scala 48:55:@3222.4]
  wire [1:0] _T_3856; // @[Bitwise.scala 48:55:@3223.4]
  wire [2:0] _T_3857; // @[Bitwise.scala 48:55:@3224.4]
  wire [3:0] _T_3858; // @[Bitwise.scala 48:55:@3225.4]
  wire [1:0] _T_3859; // @[Bitwise.scala 48:55:@3226.4]
  wire [1:0] _T_3860; // @[Bitwise.scala 48:55:@3227.4]
  wire [2:0] _T_3861; // @[Bitwise.scala 48:55:@3228.4]
  wire [1:0] _T_3862; // @[Bitwise.scala 48:55:@3229.4]
  wire [1:0] _T_3863; // @[Bitwise.scala 48:55:@3230.4]
  wire [2:0] _T_3864; // @[Bitwise.scala 48:55:@3231.4]
  wire [3:0] _T_3865; // @[Bitwise.scala 48:55:@3232.4]
  wire [4:0] _T_3866; // @[Bitwise.scala 48:55:@3233.4]
  wire [1:0] _T_3867; // @[Bitwise.scala 48:55:@3234.4]
  wire [1:0] _GEN_654; // @[Bitwise.scala 48:55:@3235.4]
  wire [2:0] _T_3868; // @[Bitwise.scala 48:55:@3235.4]
  wire [1:0] _T_3869; // @[Bitwise.scala 48:55:@3236.4]
  wire [1:0] _T_3870; // @[Bitwise.scala 48:55:@3237.4]
  wire [2:0] _T_3871; // @[Bitwise.scala 48:55:@3238.4]
  wire [3:0] _T_3872; // @[Bitwise.scala 48:55:@3239.4]
  wire [1:0] _T_3873; // @[Bitwise.scala 48:55:@3240.4]
  wire [1:0] _T_3874; // @[Bitwise.scala 48:55:@3241.4]
  wire [2:0] _T_3875; // @[Bitwise.scala 48:55:@3242.4]
  wire [1:0] _T_3876; // @[Bitwise.scala 48:55:@3243.4]
  wire [1:0] _T_3877; // @[Bitwise.scala 48:55:@3244.4]
  wire [2:0] _T_3878; // @[Bitwise.scala 48:55:@3245.4]
  wire [3:0] _T_3879; // @[Bitwise.scala 48:55:@3246.4]
  wire [4:0] _T_3880; // @[Bitwise.scala 48:55:@3247.4]
  wire [5:0] _T_3881; // @[Bitwise.scala 48:55:@3248.4]
  wire [30:0] _T_3945; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3313.4]
  wire  _T_3946; // @[Bitwise.scala 50:65:@3314.4]
  wire  _T_3947; // @[Bitwise.scala 50:65:@3315.4]
  wire  _T_3948; // @[Bitwise.scala 50:65:@3316.4]
  wire  _T_3949; // @[Bitwise.scala 50:65:@3317.4]
  wire  _T_3950; // @[Bitwise.scala 50:65:@3318.4]
  wire  _T_3951; // @[Bitwise.scala 50:65:@3319.4]
  wire  _T_3952; // @[Bitwise.scala 50:65:@3320.4]
  wire  _T_3953; // @[Bitwise.scala 50:65:@3321.4]
  wire  _T_3954; // @[Bitwise.scala 50:65:@3322.4]
  wire  _T_3955; // @[Bitwise.scala 50:65:@3323.4]
  wire  _T_3956; // @[Bitwise.scala 50:65:@3324.4]
  wire  _T_3957; // @[Bitwise.scala 50:65:@3325.4]
  wire  _T_3958; // @[Bitwise.scala 50:65:@3326.4]
  wire  _T_3959; // @[Bitwise.scala 50:65:@3327.4]
  wire  _T_3960; // @[Bitwise.scala 50:65:@3328.4]
  wire  _T_3961; // @[Bitwise.scala 50:65:@3329.4]
  wire  _T_3962; // @[Bitwise.scala 50:65:@3330.4]
  wire  _T_3963; // @[Bitwise.scala 50:65:@3331.4]
  wire  _T_3964; // @[Bitwise.scala 50:65:@3332.4]
  wire  _T_3965; // @[Bitwise.scala 50:65:@3333.4]
  wire  _T_3966; // @[Bitwise.scala 50:65:@3334.4]
  wire  _T_3967; // @[Bitwise.scala 50:65:@3335.4]
  wire  _T_3968; // @[Bitwise.scala 50:65:@3336.4]
  wire  _T_3969; // @[Bitwise.scala 50:65:@3337.4]
  wire  _T_3970; // @[Bitwise.scala 50:65:@3338.4]
  wire  _T_3971; // @[Bitwise.scala 50:65:@3339.4]
  wire  _T_3972; // @[Bitwise.scala 50:65:@3340.4]
  wire  _T_3973; // @[Bitwise.scala 50:65:@3341.4]
  wire  _T_3974; // @[Bitwise.scala 50:65:@3342.4]
  wire  _T_3975; // @[Bitwise.scala 50:65:@3343.4]
  wire  _T_3976; // @[Bitwise.scala 50:65:@3344.4]
  wire [1:0] _T_3977; // @[Bitwise.scala 48:55:@3345.4]
  wire [1:0] _GEN_655; // @[Bitwise.scala 48:55:@3346.4]
  wire [2:0] _T_3978; // @[Bitwise.scala 48:55:@3346.4]
  wire [1:0] _T_3979; // @[Bitwise.scala 48:55:@3347.4]
  wire [1:0] _T_3980; // @[Bitwise.scala 48:55:@3348.4]
  wire [2:0] _T_3981; // @[Bitwise.scala 48:55:@3349.4]
  wire [3:0] _T_3982; // @[Bitwise.scala 48:55:@3350.4]
  wire [1:0] _T_3983; // @[Bitwise.scala 48:55:@3351.4]
  wire [1:0] _T_3984; // @[Bitwise.scala 48:55:@3352.4]
  wire [2:0] _T_3985; // @[Bitwise.scala 48:55:@3353.4]
  wire [1:0] _T_3986; // @[Bitwise.scala 48:55:@3354.4]
  wire [1:0] _T_3987; // @[Bitwise.scala 48:55:@3355.4]
  wire [2:0] _T_3988; // @[Bitwise.scala 48:55:@3356.4]
  wire [3:0] _T_3989; // @[Bitwise.scala 48:55:@3357.4]
  wire [4:0] _T_3990; // @[Bitwise.scala 48:55:@3358.4]
  wire [1:0] _T_3991; // @[Bitwise.scala 48:55:@3359.4]
  wire [1:0] _T_3992; // @[Bitwise.scala 48:55:@3360.4]
  wire [2:0] _T_3993; // @[Bitwise.scala 48:55:@3361.4]
  wire [1:0] _T_3994; // @[Bitwise.scala 48:55:@3362.4]
  wire [1:0] _T_3995; // @[Bitwise.scala 48:55:@3363.4]
  wire [2:0] _T_3996; // @[Bitwise.scala 48:55:@3364.4]
  wire [3:0] _T_3997; // @[Bitwise.scala 48:55:@3365.4]
  wire [1:0] _T_3998; // @[Bitwise.scala 48:55:@3366.4]
  wire [1:0] _T_3999; // @[Bitwise.scala 48:55:@3367.4]
  wire [2:0] _T_4000; // @[Bitwise.scala 48:55:@3368.4]
  wire [1:0] _T_4001; // @[Bitwise.scala 48:55:@3369.4]
  wire [1:0] _T_4002; // @[Bitwise.scala 48:55:@3370.4]
  wire [2:0] _T_4003; // @[Bitwise.scala 48:55:@3371.4]
  wire [3:0] _T_4004; // @[Bitwise.scala 48:55:@3372.4]
  wire [4:0] _T_4005; // @[Bitwise.scala 48:55:@3373.4]
  wire [5:0] _T_4006; // @[Bitwise.scala 48:55:@3374.4]
  wire [31:0] _T_4070; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3439.4]
  wire  _T_4071; // @[Bitwise.scala 50:65:@3440.4]
  wire  _T_4072; // @[Bitwise.scala 50:65:@3441.4]
  wire  _T_4073; // @[Bitwise.scala 50:65:@3442.4]
  wire  _T_4074; // @[Bitwise.scala 50:65:@3443.4]
  wire  _T_4075; // @[Bitwise.scala 50:65:@3444.4]
  wire  _T_4076; // @[Bitwise.scala 50:65:@3445.4]
  wire  _T_4077; // @[Bitwise.scala 50:65:@3446.4]
  wire  _T_4078; // @[Bitwise.scala 50:65:@3447.4]
  wire  _T_4079; // @[Bitwise.scala 50:65:@3448.4]
  wire  _T_4080; // @[Bitwise.scala 50:65:@3449.4]
  wire  _T_4081; // @[Bitwise.scala 50:65:@3450.4]
  wire  _T_4082; // @[Bitwise.scala 50:65:@3451.4]
  wire  _T_4083; // @[Bitwise.scala 50:65:@3452.4]
  wire  _T_4084; // @[Bitwise.scala 50:65:@3453.4]
  wire  _T_4085; // @[Bitwise.scala 50:65:@3454.4]
  wire  _T_4086; // @[Bitwise.scala 50:65:@3455.4]
  wire  _T_4087; // @[Bitwise.scala 50:65:@3456.4]
  wire  _T_4088; // @[Bitwise.scala 50:65:@3457.4]
  wire  _T_4089; // @[Bitwise.scala 50:65:@3458.4]
  wire  _T_4090; // @[Bitwise.scala 50:65:@3459.4]
  wire  _T_4091; // @[Bitwise.scala 50:65:@3460.4]
  wire  _T_4092; // @[Bitwise.scala 50:65:@3461.4]
  wire  _T_4093; // @[Bitwise.scala 50:65:@3462.4]
  wire  _T_4094; // @[Bitwise.scala 50:65:@3463.4]
  wire  _T_4095; // @[Bitwise.scala 50:65:@3464.4]
  wire  _T_4096; // @[Bitwise.scala 50:65:@3465.4]
  wire  _T_4097; // @[Bitwise.scala 50:65:@3466.4]
  wire  _T_4098; // @[Bitwise.scala 50:65:@3467.4]
  wire  _T_4099; // @[Bitwise.scala 50:65:@3468.4]
  wire  _T_4100; // @[Bitwise.scala 50:65:@3469.4]
  wire  _T_4101; // @[Bitwise.scala 50:65:@3470.4]
  wire  _T_4102; // @[Bitwise.scala 50:65:@3471.4]
  wire [1:0] _T_4103; // @[Bitwise.scala 48:55:@3472.4]
  wire [1:0] _T_4104; // @[Bitwise.scala 48:55:@3473.4]
  wire [2:0] _T_4105; // @[Bitwise.scala 48:55:@3474.4]
  wire [1:0] _T_4106; // @[Bitwise.scala 48:55:@3475.4]
  wire [1:0] _T_4107; // @[Bitwise.scala 48:55:@3476.4]
  wire [2:0] _T_4108; // @[Bitwise.scala 48:55:@3477.4]
  wire [3:0] _T_4109; // @[Bitwise.scala 48:55:@3478.4]
  wire [1:0] _T_4110; // @[Bitwise.scala 48:55:@3479.4]
  wire [1:0] _T_4111; // @[Bitwise.scala 48:55:@3480.4]
  wire [2:0] _T_4112; // @[Bitwise.scala 48:55:@3481.4]
  wire [1:0] _T_4113; // @[Bitwise.scala 48:55:@3482.4]
  wire [1:0] _T_4114; // @[Bitwise.scala 48:55:@3483.4]
  wire [2:0] _T_4115; // @[Bitwise.scala 48:55:@3484.4]
  wire [3:0] _T_4116; // @[Bitwise.scala 48:55:@3485.4]
  wire [4:0] _T_4117; // @[Bitwise.scala 48:55:@3486.4]
  wire [1:0] _T_4118; // @[Bitwise.scala 48:55:@3487.4]
  wire [1:0] _T_4119; // @[Bitwise.scala 48:55:@3488.4]
  wire [2:0] _T_4120; // @[Bitwise.scala 48:55:@3489.4]
  wire [1:0] _T_4121; // @[Bitwise.scala 48:55:@3490.4]
  wire [1:0] _T_4122; // @[Bitwise.scala 48:55:@3491.4]
  wire [2:0] _T_4123; // @[Bitwise.scala 48:55:@3492.4]
  wire [3:0] _T_4124; // @[Bitwise.scala 48:55:@3493.4]
  wire [1:0] _T_4125; // @[Bitwise.scala 48:55:@3494.4]
  wire [1:0] _T_4126; // @[Bitwise.scala 48:55:@3495.4]
  wire [2:0] _T_4127; // @[Bitwise.scala 48:55:@3496.4]
  wire [1:0] _T_4128; // @[Bitwise.scala 48:55:@3497.4]
  wire [1:0] _T_4129; // @[Bitwise.scala 48:55:@3498.4]
  wire [2:0] _T_4130; // @[Bitwise.scala 48:55:@3499.4]
  wire [3:0] _T_4131; // @[Bitwise.scala 48:55:@3500.4]
  wire [4:0] _T_4132; // @[Bitwise.scala 48:55:@3501.4]
  wire [5:0] _T_4133; // @[Bitwise.scala 48:55:@3502.4]
  wire [32:0] _T_4197; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3567.4]
  wire  _T_4198; // @[Bitwise.scala 50:65:@3568.4]
  wire  _T_4199; // @[Bitwise.scala 50:65:@3569.4]
  wire  _T_4200; // @[Bitwise.scala 50:65:@3570.4]
  wire  _T_4201; // @[Bitwise.scala 50:65:@3571.4]
  wire  _T_4202; // @[Bitwise.scala 50:65:@3572.4]
  wire  _T_4203; // @[Bitwise.scala 50:65:@3573.4]
  wire  _T_4204; // @[Bitwise.scala 50:65:@3574.4]
  wire  _T_4205; // @[Bitwise.scala 50:65:@3575.4]
  wire  _T_4206; // @[Bitwise.scala 50:65:@3576.4]
  wire  _T_4207; // @[Bitwise.scala 50:65:@3577.4]
  wire  _T_4208; // @[Bitwise.scala 50:65:@3578.4]
  wire  _T_4209; // @[Bitwise.scala 50:65:@3579.4]
  wire  _T_4210; // @[Bitwise.scala 50:65:@3580.4]
  wire  _T_4211; // @[Bitwise.scala 50:65:@3581.4]
  wire  _T_4212; // @[Bitwise.scala 50:65:@3582.4]
  wire  _T_4213; // @[Bitwise.scala 50:65:@3583.4]
  wire  _T_4214; // @[Bitwise.scala 50:65:@3584.4]
  wire  _T_4215; // @[Bitwise.scala 50:65:@3585.4]
  wire  _T_4216; // @[Bitwise.scala 50:65:@3586.4]
  wire  _T_4217; // @[Bitwise.scala 50:65:@3587.4]
  wire  _T_4218; // @[Bitwise.scala 50:65:@3588.4]
  wire  _T_4219; // @[Bitwise.scala 50:65:@3589.4]
  wire  _T_4220; // @[Bitwise.scala 50:65:@3590.4]
  wire  _T_4221; // @[Bitwise.scala 50:65:@3591.4]
  wire  _T_4222; // @[Bitwise.scala 50:65:@3592.4]
  wire  _T_4223; // @[Bitwise.scala 50:65:@3593.4]
  wire  _T_4224; // @[Bitwise.scala 50:65:@3594.4]
  wire  _T_4225; // @[Bitwise.scala 50:65:@3595.4]
  wire  _T_4226; // @[Bitwise.scala 50:65:@3596.4]
  wire  _T_4227; // @[Bitwise.scala 50:65:@3597.4]
  wire  _T_4228; // @[Bitwise.scala 50:65:@3598.4]
  wire  _T_4229; // @[Bitwise.scala 50:65:@3599.4]
  wire  _T_4230; // @[Bitwise.scala 50:65:@3600.4]
  wire [1:0] _T_4231; // @[Bitwise.scala 48:55:@3601.4]
  wire [1:0] _T_4232; // @[Bitwise.scala 48:55:@3602.4]
  wire [2:0] _T_4233; // @[Bitwise.scala 48:55:@3603.4]
  wire [1:0] _T_4234; // @[Bitwise.scala 48:55:@3604.4]
  wire [1:0] _T_4235; // @[Bitwise.scala 48:55:@3605.4]
  wire [2:0] _T_4236; // @[Bitwise.scala 48:55:@3606.4]
  wire [3:0] _T_4237; // @[Bitwise.scala 48:55:@3607.4]
  wire [1:0] _T_4238; // @[Bitwise.scala 48:55:@3608.4]
  wire [1:0] _T_4239; // @[Bitwise.scala 48:55:@3609.4]
  wire [2:0] _T_4240; // @[Bitwise.scala 48:55:@3610.4]
  wire [1:0] _T_4241; // @[Bitwise.scala 48:55:@3611.4]
  wire [1:0] _T_4242; // @[Bitwise.scala 48:55:@3612.4]
  wire [2:0] _T_4243; // @[Bitwise.scala 48:55:@3613.4]
  wire [3:0] _T_4244; // @[Bitwise.scala 48:55:@3614.4]
  wire [4:0] _T_4245; // @[Bitwise.scala 48:55:@3615.4]
  wire [1:0] _T_4246; // @[Bitwise.scala 48:55:@3616.4]
  wire [1:0] _T_4247; // @[Bitwise.scala 48:55:@3617.4]
  wire [2:0] _T_4248; // @[Bitwise.scala 48:55:@3618.4]
  wire [1:0] _T_4249; // @[Bitwise.scala 48:55:@3619.4]
  wire [1:0] _T_4250; // @[Bitwise.scala 48:55:@3620.4]
  wire [2:0] _T_4251; // @[Bitwise.scala 48:55:@3621.4]
  wire [3:0] _T_4252; // @[Bitwise.scala 48:55:@3622.4]
  wire [1:0] _T_4253; // @[Bitwise.scala 48:55:@3623.4]
  wire [1:0] _T_4254; // @[Bitwise.scala 48:55:@3624.4]
  wire [2:0] _T_4255; // @[Bitwise.scala 48:55:@3625.4]
  wire [1:0] _T_4256; // @[Bitwise.scala 48:55:@3626.4]
  wire [1:0] _T_4257; // @[Bitwise.scala 48:55:@3627.4]
  wire [1:0] _GEN_656; // @[Bitwise.scala 48:55:@3628.4]
  wire [2:0] _T_4258; // @[Bitwise.scala 48:55:@3628.4]
  wire [2:0] _GEN_657; // @[Bitwise.scala 48:55:@3629.4]
  wire [3:0] _T_4259; // @[Bitwise.scala 48:55:@3629.4]
  wire [3:0] _GEN_658; // @[Bitwise.scala 48:55:@3630.4]
  wire [4:0] _T_4260; // @[Bitwise.scala 48:55:@3630.4]
  wire [4:0] _GEN_659; // @[Bitwise.scala 48:55:@3631.4]
  wire [5:0] _T_4261; // @[Bitwise.scala 48:55:@3631.4]
  wire [5:0] _GEN_660; // @[Bitwise.scala 48:55:@3632.4]
  wire [6:0] _T_4262; // @[Bitwise.scala 48:55:@3632.4]
  wire [33:0] _T_4326; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3697.4]
  wire  _T_4327; // @[Bitwise.scala 50:65:@3698.4]
  wire  _T_4328; // @[Bitwise.scala 50:65:@3699.4]
  wire  _T_4329; // @[Bitwise.scala 50:65:@3700.4]
  wire  _T_4330; // @[Bitwise.scala 50:65:@3701.4]
  wire  _T_4331; // @[Bitwise.scala 50:65:@3702.4]
  wire  _T_4332; // @[Bitwise.scala 50:65:@3703.4]
  wire  _T_4333; // @[Bitwise.scala 50:65:@3704.4]
  wire  _T_4334; // @[Bitwise.scala 50:65:@3705.4]
  wire  _T_4335; // @[Bitwise.scala 50:65:@3706.4]
  wire  _T_4336; // @[Bitwise.scala 50:65:@3707.4]
  wire  _T_4337; // @[Bitwise.scala 50:65:@3708.4]
  wire  _T_4338; // @[Bitwise.scala 50:65:@3709.4]
  wire  _T_4339; // @[Bitwise.scala 50:65:@3710.4]
  wire  _T_4340; // @[Bitwise.scala 50:65:@3711.4]
  wire  _T_4341; // @[Bitwise.scala 50:65:@3712.4]
  wire  _T_4342; // @[Bitwise.scala 50:65:@3713.4]
  wire  _T_4343; // @[Bitwise.scala 50:65:@3714.4]
  wire  _T_4344; // @[Bitwise.scala 50:65:@3715.4]
  wire  _T_4345; // @[Bitwise.scala 50:65:@3716.4]
  wire  _T_4346; // @[Bitwise.scala 50:65:@3717.4]
  wire  _T_4347; // @[Bitwise.scala 50:65:@3718.4]
  wire  _T_4348; // @[Bitwise.scala 50:65:@3719.4]
  wire  _T_4349; // @[Bitwise.scala 50:65:@3720.4]
  wire  _T_4350; // @[Bitwise.scala 50:65:@3721.4]
  wire  _T_4351; // @[Bitwise.scala 50:65:@3722.4]
  wire  _T_4352; // @[Bitwise.scala 50:65:@3723.4]
  wire  _T_4353; // @[Bitwise.scala 50:65:@3724.4]
  wire  _T_4354; // @[Bitwise.scala 50:65:@3725.4]
  wire  _T_4355; // @[Bitwise.scala 50:65:@3726.4]
  wire  _T_4356; // @[Bitwise.scala 50:65:@3727.4]
  wire  _T_4357; // @[Bitwise.scala 50:65:@3728.4]
  wire  _T_4358; // @[Bitwise.scala 50:65:@3729.4]
  wire  _T_4359; // @[Bitwise.scala 50:65:@3730.4]
  wire  _T_4360; // @[Bitwise.scala 50:65:@3731.4]
  wire [1:0] _T_4361; // @[Bitwise.scala 48:55:@3732.4]
  wire [1:0] _T_4362; // @[Bitwise.scala 48:55:@3733.4]
  wire [2:0] _T_4363; // @[Bitwise.scala 48:55:@3734.4]
  wire [1:0] _T_4364; // @[Bitwise.scala 48:55:@3735.4]
  wire [1:0] _T_4365; // @[Bitwise.scala 48:55:@3736.4]
  wire [2:0] _T_4366; // @[Bitwise.scala 48:55:@3737.4]
  wire [3:0] _T_4367; // @[Bitwise.scala 48:55:@3738.4]
  wire [1:0] _T_4368; // @[Bitwise.scala 48:55:@3739.4]
  wire [1:0] _T_4369; // @[Bitwise.scala 48:55:@3740.4]
  wire [2:0] _T_4370; // @[Bitwise.scala 48:55:@3741.4]
  wire [1:0] _T_4371; // @[Bitwise.scala 48:55:@3742.4]
  wire [1:0] _T_4372; // @[Bitwise.scala 48:55:@3743.4]
  wire [1:0] _GEN_661; // @[Bitwise.scala 48:55:@3744.4]
  wire [2:0] _T_4373; // @[Bitwise.scala 48:55:@3744.4]
  wire [2:0] _GEN_662; // @[Bitwise.scala 48:55:@3745.4]
  wire [3:0] _T_4374; // @[Bitwise.scala 48:55:@3745.4]
  wire [3:0] _GEN_663; // @[Bitwise.scala 48:55:@3746.4]
  wire [4:0] _T_4375; // @[Bitwise.scala 48:55:@3746.4]
  wire [4:0] _GEN_664; // @[Bitwise.scala 48:55:@3747.4]
  wire [5:0] _T_4376; // @[Bitwise.scala 48:55:@3747.4]
  wire [1:0] _T_4377; // @[Bitwise.scala 48:55:@3748.4]
  wire [1:0] _T_4378; // @[Bitwise.scala 48:55:@3749.4]
  wire [2:0] _T_4379; // @[Bitwise.scala 48:55:@3750.4]
  wire [1:0] _T_4380; // @[Bitwise.scala 48:55:@3751.4]
  wire [1:0] _T_4381; // @[Bitwise.scala 48:55:@3752.4]
  wire [2:0] _T_4382; // @[Bitwise.scala 48:55:@3753.4]
  wire [3:0] _T_4383; // @[Bitwise.scala 48:55:@3754.4]
  wire [1:0] _T_4384; // @[Bitwise.scala 48:55:@3755.4]
  wire [1:0] _T_4385; // @[Bitwise.scala 48:55:@3756.4]
  wire [2:0] _T_4386; // @[Bitwise.scala 48:55:@3757.4]
  wire [1:0] _T_4387; // @[Bitwise.scala 48:55:@3758.4]
  wire [1:0] _T_4388; // @[Bitwise.scala 48:55:@3759.4]
  wire [1:0] _GEN_665; // @[Bitwise.scala 48:55:@3760.4]
  wire [2:0] _T_4389; // @[Bitwise.scala 48:55:@3760.4]
  wire [2:0] _GEN_666; // @[Bitwise.scala 48:55:@3761.4]
  wire [3:0] _T_4390; // @[Bitwise.scala 48:55:@3761.4]
  wire [3:0] _GEN_667; // @[Bitwise.scala 48:55:@3762.4]
  wire [4:0] _T_4391; // @[Bitwise.scala 48:55:@3762.4]
  wire [4:0] _GEN_668; // @[Bitwise.scala 48:55:@3763.4]
  wire [5:0] _T_4392; // @[Bitwise.scala 48:55:@3763.4]
  wire [6:0] _T_4393; // @[Bitwise.scala 48:55:@3764.4]
  wire [34:0] _T_4457; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3829.4]
  wire  _T_4458; // @[Bitwise.scala 50:65:@3830.4]
  wire  _T_4459; // @[Bitwise.scala 50:65:@3831.4]
  wire  _T_4460; // @[Bitwise.scala 50:65:@3832.4]
  wire  _T_4461; // @[Bitwise.scala 50:65:@3833.4]
  wire  _T_4462; // @[Bitwise.scala 50:65:@3834.4]
  wire  _T_4463; // @[Bitwise.scala 50:65:@3835.4]
  wire  _T_4464; // @[Bitwise.scala 50:65:@3836.4]
  wire  _T_4465; // @[Bitwise.scala 50:65:@3837.4]
  wire  _T_4466; // @[Bitwise.scala 50:65:@3838.4]
  wire  _T_4467; // @[Bitwise.scala 50:65:@3839.4]
  wire  _T_4468; // @[Bitwise.scala 50:65:@3840.4]
  wire  _T_4469; // @[Bitwise.scala 50:65:@3841.4]
  wire  _T_4470; // @[Bitwise.scala 50:65:@3842.4]
  wire  _T_4471; // @[Bitwise.scala 50:65:@3843.4]
  wire  _T_4472; // @[Bitwise.scala 50:65:@3844.4]
  wire  _T_4473; // @[Bitwise.scala 50:65:@3845.4]
  wire  _T_4474; // @[Bitwise.scala 50:65:@3846.4]
  wire  _T_4475; // @[Bitwise.scala 50:65:@3847.4]
  wire  _T_4476; // @[Bitwise.scala 50:65:@3848.4]
  wire  _T_4477; // @[Bitwise.scala 50:65:@3849.4]
  wire  _T_4478; // @[Bitwise.scala 50:65:@3850.4]
  wire  _T_4479; // @[Bitwise.scala 50:65:@3851.4]
  wire  _T_4480; // @[Bitwise.scala 50:65:@3852.4]
  wire  _T_4481; // @[Bitwise.scala 50:65:@3853.4]
  wire  _T_4482; // @[Bitwise.scala 50:65:@3854.4]
  wire  _T_4483; // @[Bitwise.scala 50:65:@3855.4]
  wire  _T_4484; // @[Bitwise.scala 50:65:@3856.4]
  wire  _T_4485; // @[Bitwise.scala 50:65:@3857.4]
  wire  _T_4486; // @[Bitwise.scala 50:65:@3858.4]
  wire  _T_4487; // @[Bitwise.scala 50:65:@3859.4]
  wire  _T_4488; // @[Bitwise.scala 50:65:@3860.4]
  wire  _T_4489; // @[Bitwise.scala 50:65:@3861.4]
  wire  _T_4490; // @[Bitwise.scala 50:65:@3862.4]
  wire  _T_4491; // @[Bitwise.scala 50:65:@3863.4]
  wire  _T_4492; // @[Bitwise.scala 50:65:@3864.4]
  wire [1:0] _T_4493; // @[Bitwise.scala 48:55:@3865.4]
  wire [1:0] _T_4494; // @[Bitwise.scala 48:55:@3866.4]
  wire [2:0] _T_4495; // @[Bitwise.scala 48:55:@3867.4]
  wire [1:0] _T_4496; // @[Bitwise.scala 48:55:@3868.4]
  wire [1:0] _T_4497; // @[Bitwise.scala 48:55:@3869.4]
  wire [2:0] _T_4498; // @[Bitwise.scala 48:55:@3870.4]
  wire [3:0] _T_4499; // @[Bitwise.scala 48:55:@3871.4]
  wire [1:0] _T_4500; // @[Bitwise.scala 48:55:@3872.4]
  wire [1:0] _T_4501; // @[Bitwise.scala 48:55:@3873.4]
  wire [2:0] _T_4502; // @[Bitwise.scala 48:55:@3874.4]
  wire [1:0] _T_4503; // @[Bitwise.scala 48:55:@3875.4]
  wire [1:0] _T_4504; // @[Bitwise.scala 48:55:@3876.4]
  wire [1:0] _GEN_669; // @[Bitwise.scala 48:55:@3877.4]
  wire [2:0] _T_4505; // @[Bitwise.scala 48:55:@3877.4]
  wire [2:0] _GEN_670; // @[Bitwise.scala 48:55:@3878.4]
  wire [3:0] _T_4506; // @[Bitwise.scala 48:55:@3878.4]
  wire [3:0] _GEN_671; // @[Bitwise.scala 48:55:@3879.4]
  wire [4:0] _T_4507; // @[Bitwise.scala 48:55:@3879.4]
  wire [4:0] _GEN_672; // @[Bitwise.scala 48:55:@3880.4]
  wire [5:0] _T_4508; // @[Bitwise.scala 48:55:@3880.4]
  wire [1:0] _T_4509; // @[Bitwise.scala 48:55:@3881.4]
  wire [1:0] _T_4510; // @[Bitwise.scala 48:55:@3882.4]
  wire [2:0] _T_4511; // @[Bitwise.scala 48:55:@3883.4]
  wire [1:0] _T_4512; // @[Bitwise.scala 48:55:@3884.4]
  wire [1:0] _T_4513; // @[Bitwise.scala 48:55:@3885.4]
  wire [1:0] _GEN_673; // @[Bitwise.scala 48:55:@3886.4]
  wire [2:0] _T_4514; // @[Bitwise.scala 48:55:@3886.4]
  wire [2:0] _GEN_674; // @[Bitwise.scala 48:55:@3887.4]
  wire [3:0] _T_4515; // @[Bitwise.scala 48:55:@3887.4]
  wire [3:0] _GEN_675; // @[Bitwise.scala 48:55:@3888.4]
  wire [4:0] _T_4516; // @[Bitwise.scala 48:55:@3888.4]
  wire [1:0] _T_4517; // @[Bitwise.scala 48:55:@3889.4]
  wire [1:0] _T_4518; // @[Bitwise.scala 48:55:@3890.4]
  wire [2:0] _T_4519; // @[Bitwise.scala 48:55:@3891.4]
  wire [1:0] _T_4520; // @[Bitwise.scala 48:55:@3892.4]
  wire [1:0] _T_4521; // @[Bitwise.scala 48:55:@3893.4]
  wire [1:0] _GEN_676; // @[Bitwise.scala 48:55:@3894.4]
  wire [2:0] _T_4522; // @[Bitwise.scala 48:55:@3894.4]
  wire [2:0] _GEN_677; // @[Bitwise.scala 48:55:@3895.4]
  wire [3:0] _T_4523; // @[Bitwise.scala 48:55:@3895.4]
  wire [3:0] _GEN_678; // @[Bitwise.scala 48:55:@3896.4]
  wire [4:0] _T_4524; // @[Bitwise.scala 48:55:@3896.4]
  wire [5:0] _T_4525; // @[Bitwise.scala 48:55:@3897.4]
  wire [6:0] _T_4526; // @[Bitwise.scala 48:55:@3898.4]
  wire [35:0] _T_4590; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3963.4]
  wire  _T_4591; // @[Bitwise.scala 50:65:@3964.4]
  wire  _T_4592; // @[Bitwise.scala 50:65:@3965.4]
  wire  _T_4593; // @[Bitwise.scala 50:65:@3966.4]
  wire  _T_4594; // @[Bitwise.scala 50:65:@3967.4]
  wire  _T_4595; // @[Bitwise.scala 50:65:@3968.4]
  wire  _T_4596; // @[Bitwise.scala 50:65:@3969.4]
  wire  _T_4597; // @[Bitwise.scala 50:65:@3970.4]
  wire  _T_4598; // @[Bitwise.scala 50:65:@3971.4]
  wire  _T_4599; // @[Bitwise.scala 50:65:@3972.4]
  wire  _T_4600; // @[Bitwise.scala 50:65:@3973.4]
  wire  _T_4601; // @[Bitwise.scala 50:65:@3974.4]
  wire  _T_4602; // @[Bitwise.scala 50:65:@3975.4]
  wire  _T_4603; // @[Bitwise.scala 50:65:@3976.4]
  wire  _T_4604; // @[Bitwise.scala 50:65:@3977.4]
  wire  _T_4605; // @[Bitwise.scala 50:65:@3978.4]
  wire  _T_4606; // @[Bitwise.scala 50:65:@3979.4]
  wire  _T_4607; // @[Bitwise.scala 50:65:@3980.4]
  wire  _T_4608; // @[Bitwise.scala 50:65:@3981.4]
  wire  _T_4609; // @[Bitwise.scala 50:65:@3982.4]
  wire  _T_4610; // @[Bitwise.scala 50:65:@3983.4]
  wire  _T_4611; // @[Bitwise.scala 50:65:@3984.4]
  wire  _T_4612; // @[Bitwise.scala 50:65:@3985.4]
  wire  _T_4613; // @[Bitwise.scala 50:65:@3986.4]
  wire  _T_4614; // @[Bitwise.scala 50:65:@3987.4]
  wire  _T_4615; // @[Bitwise.scala 50:65:@3988.4]
  wire  _T_4616; // @[Bitwise.scala 50:65:@3989.4]
  wire  _T_4617; // @[Bitwise.scala 50:65:@3990.4]
  wire  _T_4618; // @[Bitwise.scala 50:65:@3991.4]
  wire  _T_4619; // @[Bitwise.scala 50:65:@3992.4]
  wire  _T_4620; // @[Bitwise.scala 50:65:@3993.4]
  wire  _T_4621; // @[Bitwise.scala 50:65:@3994.4]
  wire  _T_4622; // @[Bitwise.scala 50:65:@3995.4]
  wire  _T_4623; // @[Bitwise.scala 50:65:@3996.4]
  wire  _T_4624; // @[Bitwise.scala 50:65:@3997.4]
  wire  _T_4625; // @[Bitwise.scala 50:65:@3998.4]
  wire  _T_4626; // @[Bitwise.scala 50:65:@3999.4]
  wire [1:0] _T_4627; // @[Bitwise.scala 48:55:@4000.4]
  wire [1:0] _T_4628; // @[Bitwise.scala 48:55:@4001.4]
  wire [2:0] _T_4629; // @[Bitwise.scala 48:55:@4002.4]
  wire [1:0] _T_4630; // @[Bitwise.scala 48:55:@4003.4]
  wire [1:0] _T_4631; // @[Bitwise.scala 48:55:@4004.4]
  wire [1:0] _GEN_679; // @[Bitwise.scala 48:55:@4005.4]
  wire [2:0] _T_4632; // @[Bitwise.scala 48:55:@4005.4]
  wire [2:0] _GEN_680; // @[Bitwise.scala 48:55:@4006.4]
  wire [3:0] _T_4633; // @[Bitwise.scala 48:55:@4006.4]
  wire [3:0] _GEN_681; // @[Bitwise.scala 48:55:@4007.4]
  wire [4:0] _T_4634; // @[Bitwise.scala 48:55:@4007.4]
  wire [1:0] _T_4635; // @[Bitwise.scala 48:55:@4008.4]
  wire [1:0] _T_4636; // @[Bitwise.scala 48:55:@4009.4]
  wire [2:0] _T_4637; // @[Bitwise.scala 48:55:@4010.4]
  wire [1:0] _T_4638; // @[Bitwise.scala 48:55:@4011.4]
  wire [1:0] _T_4639; // @[Bitwise.scala 48:55:@4012.4]
  wire [1:0] _GEN_682; // @[Bitwise.scala 48:55:@4013.4]
  wire [2:0] _T_4640; // @[Bitwise.scala 48:55:@4013.4]
  wire [2:0] _GEN_683; // @[Bitwise.scala 48:55:@4014.4]
  wire [3:0] _T_4641; // @[Bitwise.scala 48:55:@4014.4]
  wire [3:0] _GEN_684; // @[Bitwise.scala 48:55:@4015.4]
  wire [4:0] _T_4642; // @[Bitwise.scala 48:55:@4015.4]
  wire [5:0] _T_4643; // @[Bitwise.scala 48:55:@4016.4]
  wire [1:0] _T_4644; // @[Bitwise.scala 48:55:@4017.4]
  wire [1:0] _T_4645; // @[Bitwise.scala 48:55:@4018.4]
  wire [2:0] _T_4646; // @[Bitwise.scala 48:55:@4019.4]
  wire [1:0] _T_4647; // @[Bitwise.scala 48:55:@4020.4]
  wire [1:0] _T_4648; // @[Bitwise.scala 48:55:@4021.4]
  wire [1:0] _GEN_685; // @[Bitwise.scala 48:55:@4022.4]
  wire [2:0] _T_4649; // @[Bitwise.scala 48:55:@4022.4]
  wire [2:0] _GEN_686; // @[Bitwise.scala 48:55:@4023.4]
  wire [3:0] _T_4650; // @[Bitwise.scala 48:55:@4023.4]
  wire [3:0] _GEN_687; // @[Bitwise.scala 48:55:@4024.4]
  wire [4:0] _T_4651; // @[Bitwise.scala 48:55:@4024.4]
  wire [1:0] _T_4652; // @[Bitwise.scala 48:55:@4025.4]
  wire [1:0] _T_4653; // @[Bitwise.scala 48:55:@4026.4]
  wire [2:0] _T_4654; // @[Bitwise.scala 48:55:@4027.4]
  wire [1:0] _T_4655; // @[Bitwise.scala 48:55:@4028.4]
  wire [1:0] _T_4656; // @[Bitwise.scala 48:55:@4029.4]
  wire [1:0] _GEN_688; // @[Bitwise.scala 48:55:@4030.4]
  wire [2:0] _T_4657; // @[Bitwise.scala 48:55:@4030.4]
  wire [2:0] _GEN_689; // @[Bitwise.scala 48:55:@4031.4]
  wire [3:0] _T_4658; // @[Bitwise.scala 48:55:@4031.4]
  wire [3:0] _GEN_690; // @[Bitwise.scala 48:55:@4032.4]
  wire [4:0] _T_4659; // @[Bitwise.scala 48:55:@4032.4]
  wire [5:0] _T_4660; // @[Bitwise.scala 48:55:@4033.4]
  wire [6:0] _T_4661; // @[Bitwise.scala 48:55:@4034.4]
  wire [36:0] _T_4725; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4099.4]
  wire  _T_4726; // @[Bitwise.scala 50:65:@4100.4]
  wire  _T_4727; // @[Bitwise.scala 50:65:@4101.4]
  wire  _T_4728; // @[Bitwise.scala 50:65:@4102.4]
  wire  _T_4729; // @[Bitwise.scala 50:65:@4103.4]
  wire  _T_4730; // @[Bitwise.scala 50:65:@4104.4]
  wire  _T_4731; // @[Bitwise.scala 50:65:@4105.4]
  wire  _T_4732; // @[Bitwise.scala 50:65:@4106.4]
  wire  _T_4733; // @[Bitwise.scala 50:65:@4107.4]
  wire  _T_4734; // @[Bitwise.scala 50:65:@4108.4]
  wire  _T_4735; // @[Bitwise.scala 50:65:@4109.4]
  wire  _T_4736; // @[Bitwise.scala 50:65:@4110.4]
  wire  _T_4737; // @[Bitwise.scala 50:65:@4111.4]
  wire  _T_4738; // @[Bitwise.scala 50:65:@4112.4]
  wire  _T_4739; // @[Bitwise.scala 50:65:@4113.4]
  wire  _T_4740; // @[Bitwise.scala 50:65:@4114.4]
  wire  _T_4741; // @[Bitwise.scala 50:65:@4115.4]
  wire  _T_4742; // @[Bitwise.scala 50:65:@4116.4]
  wire  _T_4743; // @[Bitwise.scala 50:65:@4117.4]
  wire  _T_4744; // @[Bitwise.scala 50:65:@4118.4]
  wire  _T_4745; // @[Bitwise.scala 50:65:@4119.4]
  wire  _T_4746; // @[Bitwise.scala 50:65:@4120.4]
  wire  _T_4747; // @[Bitwise.scala 50:65:@4121.4]
  wire  _T_4748; // @[Bitwise.scala 50:65:@4122.4]
  wire  _T_4749; // @[Bitwise.scala 50:65:@4123.4]
  wire  _T_4750; // @[Bitwise.scala 50:65:@4124.4]
  wire  _T_4751; // @[Bitwise.scala 50:65:@4125.4]
  wire  _T_4752; // @[Bitwise.scala 50:65:@4126.4]
  wire  _T_4753; // @[Bitwise.scala 50:65:@4127.4]
  wire  _T_4754; // @[Bitwise.scala 50:65:@4128.4]
  wire  _T_4755; // @[Bitwise.scala 50:65:@4129.4]
  wire  _T_4756; // @[Bitwise.scala 50:65:@4130.4]
  wire  _T_4757; // @[Bitwise.scala 50:65:@4131.4]
  wire  _T_4758; // @[Bitwise.scala 50:65:@4132.4]
  wire  _T_4759; // @[Bitwise.scala 50:65:@4133.4]
  wire  _T_4760; // @[Bitwise.scala 50:65:@4134.4]
  wire  _T_4761; // @[Bitwise.scala 50:65:@4135.4]
  wire  _T_4762; // @[Bitwise.scala 50:65:@4136.4]
  wire [1:0] _T_4763; // @[Bitwise.scala 48:55:@4137.4]
  wire [1:0] _T_4764; // @[Bitwise.scala 48:55:@4138.4]
  wire [2:0] _T_4765; // @[Bitwise.scala 48:55:@4139.4]
  wire [1:0] _T_4766; // @[Bitwise.scala 48:55:@4140.4]
  wire [1:0] _T_4767; // @[Bitwise.scala 48:55:@4141.4]
  wire [1:0] _GEN_691; // @[Bitwise.scala 48:55:@4142.4]
  wire [2:0] _T_4768; // @[Bitwise.scala 48:55:@4142.4]
  wire [2:0] _GEN_692; // @[Bitwise.scala 48:55:@4143.4]
  wire [3:0] _T_4769; // @[Bitwise.scala 48:55:@4143.4]
  wire [3:0] _GEN_693; // @[Bitwise.scala 48:55:@4144.4]
  wire [4:0] _T_4770; // @[Bitwise.scala 48:55:@4144.4]
  wire [1:0] _T_4771; // @[Bitwise.scala 48:55:@4145.4]
  wire [1:0] _T_4772; // @[Bitwise.scala 48:55:@4146.4]
  wire [2:0] _T_4773; // @[Bitwise.scala 48:55:@4147.4]
  wire [1:0] _T_4774; // @[Bitwise.scala 48:55:@4148.4]
  wire [1:0] _T_4775; // @[Bitwise.scala 48:55:@4149.4]
  wire [1:0] _GEN_694; // @[Bitwise.scala 48:55:@4150.4]
  wire [2:0] _T_4776; // @[Bitwise.scala 48:55:@4150.4]
  wire [2:0] _GEN_695; // @[Bitwise.scala 48:55:@4151.4]
  wire [3:0] _T_4777; // @[Bitwise.scala 48:55:@4151.4]
  wire [3:0] _GEN_696; // @[Bitwise.scala 48:55:@4152.4]
  wire [4:0] _T_4778; // @[Bitwise.scala 48:55:@4152.4]
  wire [5:0] _T_4779; // @[Bitwise.scala 48:55:@4153.4]
  wire [1:0] _T_4780; // @[Bitwise.scala 48:55:@4154.4]
  wire [1:0] _T_4781; // @[Bitwise.scala 48:55:@4155.4]
  wire [2:0] _T_4782; // @[Bitwise.scala 48:55:@4156.4]
  wire [1:0] _T_4783; // @[Bitwise.scala 48:55:@4157.4]
  wire [1:0] _T_4784; // @[Bitwise.scala 48:55:@4158.4]
  wire [1:0] _GEN_697; // @[Bitwise.scala 48:55:@4159.4]
  wire [2:0] _T_4785; // @[Bitwise.scala 48:55:@4159.4]
  wire [2:0] _GEN_698; // @[Bitwise.scala 48:55:@4160.4]
  wire [3:0] _T_4786; // @[Bitwise.scala 48:55:@4160.4]
  wire [3:0] _GEN_699; // @[Bitwise.scala 48:55:@4161.4]
  wire [4:0] _T_4787; // @[Bitwise.scala 48:55:@4161.4]
  wire [1:0] _T_4788; // @[Bitwise.scala 48:55:@4162.4]
  wire [1:0] _T_4789; // @[Bitwise.scala 48:55:@4163.4]
  wire [1:0] _GEN_700; // @[Bitwise.scala 48:55:@4164.4]
  wire [2:0] _T_4790; // @[Bitwise.scala 48:55:@4164.4]
  wire [2:0] _GEN_701; // @[Bitwise.scala 48:55:@4165.4]
  wire [3:0] _T_4791; // @[Bitwise.scala 48:55:@4165.4]
  wire [1:0] _T_4792; // @[Bitwise.scala 48:55:@4166.4]
  wire [1:0] _T_4793; // @[Bitwise.scala 48:55:@4167.4]
  wire [1:0] _GEN_702; // @[Bitwise.scala 48:55:@4168.4]
  wire [2:0] _T_4794; // @[Bitwise.scala 48:55:@4168.4]
  wire [2:0] _GEN_703; // @[Bitwise.scala 48:55:@4169.4]
  wire [3:0] _T_4795; // @[Bitwise.scala 48:55:@4169.4]
  wire [4:0] _T_4796; // @[Bitwise.scala 48:55:@4170.4]
  wire [5:0] _T_4797; // @[Bitwise.scala 48:55:@4171.4]
  wire [6:0] _T_4798; // @[Bitwise.scala 48:55:@4172.4]
  wire [37:0] _T_4862; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4237.4]
  wire  _T_4863; // @[Bitwise.scala 50:65:@4238.4]
  wire  _T_4864; // @[Bitwise.scala 50:65:@4239.4]
  wire  _T_4865; // @[Bitwise.scala 50:65:@4240.4]
  wire  _T_4866; // @[Bitwise.scala 50:65:@4241.4]
  wire  _T_4867; // @[Bitwise.scala 50:65:@4242.4]
  wire  _T_4868; // @[Bitwise.scala 50:65:@4243.4]
  wire  _T_4869; // @[Bitwise.scala 50:65:@4244.4]
  wire  _T_4870; // @[Bitwise.scala 50:65:@4245.4]
  wire  _T_4871; // @[Bitwise.scala 50:65:@4246.4]
  wire  _T_4872; // @[Bitwise.scala 50:65:@4247.4]
  wire  _T_4873; // @[Bitwise.scala 50:65:@4248.4]
  wire  _T_4874; // @[Bitwise.scala 50:65:@4249.4]
  wire  _T_4875; // @[Bitwise.scala 50:65:@4250.4]
  wire  _T_4876; // @[Bitwise.scala 50:65:@4251.4]
  wire  _T_4877; // @[Bitwise.scala 50:65:@4252.4]
  wire  _T_4878; // @[Bitwise.scala 50:65:@4253.4]
  wire  _T_4879; // @[Bitwise.scala 50:65:@4254.4]
  wire  _T_4880; // @[Bitwise.scala 50:65:@4255.4]
  wire  _T_4881; // @[Bitwise.scala 50:65:@4256.4]
  wire  _T_4882; // @[Bitwise.scala 50:65:@4257.4]
  wire  _T_4883; // @[Bitwise.scala 50:65:@4258.4]
  wire  _T_4884; // @[Bitwise.scala 50:65:@4259.4]
  wire  _T_4885; // @[Bitwise.scala 50:65:@4260.4]
  wire  _T_4886; // @[Bitwise.scala 50:65:@4261.4]
  wire  _T_4887; // @[Bitwise.scala 50:65:@4262.4]
  wire  _T_4888; // @[Bitwise.scala 50:65:@4263.4]
  wire  _T_4889; // @[Bitwise.scala 50:65:@4264.4]
  wire  _T_4890; // @[Bitwise.scala 50:65:@4265.4]
  wire  _T_4891; // @[Bitwise.scala 50:65:@4266.4]
  wire  _T_4892; // @[Bitwise.scala 50:65:@4267.4]
  wire  _T_4893; // @[Bitwise.scala 50:65:@4268.4]
  wire  _T_4894; // @[Bitwise.scala 50:65:@4269.4]
  wire  _T_4895; // @[Bitwise.scala 50:65:@4270.4]
  wire  _T_4896; // @[Bitwise.scala 50:65:@4271.4]
  wire  _T_4897; // @[Bitwise.scala 50:65:@4272.4]
  wire  _T_4898; // @[Bitwise.scala 50:65:@4273.4]
  wire  _T_4899; // @[Bitwise.scala 50:65:@4274.4]
  wire  _T_4900; // @[Bitwise.scala 50:65:@4275.4]
  wire [1:0] _T_4901; // @[Bitwise.scala 48:55:@4276.4]
  wire [1:0] _T_4902; // @[Bitwise.scala 48:55:@4277.4]
  wire [2:0] _T_4903; // @[Bitwise.scala 48:55:@4278.4]
  wire [1:0] _T_4904; // @[Bitwise.scala 48:55:@4279.4]
  wire [1:0] _T_4905; // @[Bitwise.scala 48:55:@4280.4]
  wire [1:0] _GEN_704; // @[Bitwise.scala 48:55:@4281.4]
  wire [2:0] _T_4906; // @[Bitwise.scala 48:55:@4281.4]
  wire [2:0] _GEN_705; // @[Bitwise.scala 48:55:@4282.4]
  wire [3:0] _T_4907; // @[Bitwise.scala 48:55:@4282.4]
  wire [3:0] _GEN_706; // @[Bitwise.scala 48:55:@4283.4]
  wire [4:0] _T_4908; // @[Bitwise.scala 48:55:@4283.4]
  wire [1:0] _T_4909; // @[Bitwise.scala 48:55:@4284.4]
  wire [1:0] _T_4910; // @[Bitwise.scala 48:55:@4285.4]
  wire [1:0] _GEN_707; // @[Bitwise.scala 48:55:@4286.4]
  wire [2:0] _T_4911; // @[Bitwise.scala 48:55:@4286.4]
  wire [2:0] _GEN_708; // @[Bitwise.scala 48:55:@4287.4]
  wire [3:0] _T_4912; // @[Bitwise.scala 48:55:@4287.4]
  wire [1:0] _T_4913; // @[Bitwise.scala 48:55:@4288.4]
  wire [1:0] _T_4914; // @[Bitwise.scala 48:55:@4289.4]
  wire [1:0] _GEN_709; // @[Bitwise.scala 48:55:@4290.4]
  wire [2:0] _T_4915; // @[Bitwise.scala 48:55:@4290.4]
  wire [2:0] _GEN_710; // @[Bitwise.scala 48:55:@4291.4]
  wire [3:0] _T_4916; // @[Bitwise.scala 48:55:@4291.4]
  wire [4:0] _T_4917; // @[Bitwise.scala 48:55:@4292.4]
  wire [5:0] _T_4918; // @[Bitwise.scala 48:55:@4293.4]
  wire [1:0] _T_4919; // @[Bitwise.scala 48:55:@4294.4]
  wire [1:0] _T_4920; // @[Bitwise.scala 48:55:@4295.4]
  wire [2:0] _T_4921; // @[Bitwise.scala 48:55:@4296.4]
  wire [1:0] _T_4922; // @[Bitwise.scala 48:55:@4297.4]
  wire [1:0] _T_4923; // @[Bitwise.scala 48:55:@4298.4]
  wire [1:0] _GEN_711; // @[Bitwise.scala 48:55:@4299.4]
  wire [2:0] _T_4924; // @[Bitwise.scala 48:55:@4299.4]
  wire [2:0] _GEN_712; // @[Bitwise.scala 48:55:@4300.4]
  wire [3:0] _T_4925; // @[Bitwise.scala 48:55:@4300.4]
  wire [3:0] _GEN_713; // @[Bitwise.scala 48:55:@4301.4]
  wire [4:0] _T_4926; // @[Bitwise.scala 48:55:@4301.4]
  wire [1:0] _T_4927; // @[Bitwise.scala 48:55:@4302.4]
  wire [1:0] _T_4928; // @[Bitwise.scala 48:55:@4303.4]
  wire [1:0] _GEN_714; // @[Bitwise.scala 48:55:@4304.4]
  wire [2:0] _T_4929; // @[Bitwise.scala 48:55:@4304.4]
  wire [2:0] _GEN_715; // @[Bitwise.scala 48:55:@4305.4]
  wire [3:0] _T_4930; // @[Bitwise.scala 48:55:@4305.4]
  wire [1:0] _T_4931; // @[Bitwise.scala 48:55:@4306.4]
  wire [1:0] _T_4932; // @[Bitwise.scala 48:55:@4307.4]
  wire [1:0] _GEN_716; // @[Bitwise.scala 48:55:@4308.4]
  wire [2:0] _T_4933; // @[Bitwise.scala 48:55:@4308.4]
  wire [2:0] _GEN_717; // @[Bitwise.scala 48:55:@4309.4]
  wire [3:0] _T_4934; // @[Bitwise.scala 48:55:@4309.4]
  wire [4:0] _T_4935; // @[Bitwise.scala 48:55:@4310.4]
  wire [5:0] _T_4936; // @[Bitwise.scala 48:55:@4311.4]
  wire [6:0] _T_4937; // @[Bitwise.scala 48:55:@4312.4]
  wire [38:0] _T_5001; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4377.4]
  wire  _T_5002; // @[Bitwise.scala 50:65:@4378.4]
  wire  _T_5003; // @[Bitwise.scala 50:65:@4379.4]
  wire  _T_5004; // @[Bitwise.scala 50:65:@4380.4]
  wire  _T_5005; // @[Bitwise.scala 50:65:@4381.4]
  wire  _T_5006; // @[Bitwise.scala 50:65:@4382.4]
  wire  _T_5007; // @[Bitwise.scala 50:65:@4383.4]
  wire  _T_5008; // @[Bitwise.scala 50:65:@4384.4]
  wire  _T_5009; // @[Bitwise.scala 50:65:@4385.4]
  wire  _T_5010; // @[Bitwise.scala 50:65:@4386.4]
  wire  _T_5011; // @[Bitwise.scala 50:65:@4387.4]
  wire  _T_5012; // @[Bitwise.scala 50:65:@4388.4]
  wire  _T_5013; // @[Bitwise.scala 50:65:@4389.4]
  wire  _T_5014; // @[Bitwise.scala 50:65:@4390.4]
  wire  _T_5015; // @[Bitwise.scala 50:65:@4391.4]
  wire  _T_5016; // @[Bitwise.scala 50:65:@4392.4]
  wire  _T_5017; // @[Bitwise.scala 50:65:@4393.4]
  wire  _T_5018; // @[Bitwise.scala 50:65:@4394.4]
  wire  _T_5019; // @[Bitwise.scala 50:65:@4395.4]
  wire  _T_5020; // @[Bitwise.scala 50:65:@4396.4]
  wire  _T_5021; // @[Bitwise.scala 50:65:@4397.4]
  wire  _T_5022; // @[Bitwise.scala 50:65:@4398.4]
  wire  _T_5023; // @[Bitwise.scala 50:65:@4399.4]
  wire  _T_5024; // @[Bitwise.scala 50:65:@4400.4]
  wire  _T_5025; // @[Bitwise.scala 50:65:@4401.4]
  wire  _T_5026; // @[Bitwise.scala 50:65:@4402.4]
  wire  _T_5027; // @[Bitwise.scala 50:65:@4403.4]
  wire  _T_5028; // @[Bitwise.scala 50:65:@4404.4]
  wire  _T_5029; // @[Bitwise.scala 50:65:@4405.4]
  wire  _T_5030; // @[Bitwise.scala 50:65:@4406.4]
  wire  _T_5031; // @[Bitwise.scala 50:65:@4407.4]
  wire  _T_5032; // @[Bitwise.scala 50:65:@4408.4]
  wire  _T_5033; // @[Bitwise.scala 50:65:@4409.4]
  wire  _T_5034; // @[Bitwise.scala 50:65:@4410.4]
  wire  _T_5035; // @[Bitwise.scala 50:65:@4411.4]
  wire  _T_5036; // @[Bitwise.scala 50:65:@4412.4]
  wire  _T_5037; // @[Bitwise.scala 50:65:@4413.4]
  wire  _T_5038; // @[Bitwise.scala 50:65:@4414.4]
  wire  _T_5039; // @[Bitwise.scala 50:65:@4415.4]
  wire  _T_5040; // @[Bitwise.scala 50:65:@4416.4]
  wire [1:0] _T_5041; // @[Bitwise.scala 48:55:@4417.4]
  wire [1:0] _T_5042; // @[Bitwise.scala 48:55:@4418.4]
  wire [2:0] _T_5043; // @[Bitwise.scala 48:55:@4419.4]
  wire [1:0] _T_5044; // @[Bitwise.scala 48:55:@4420.4]
  wire [1:0] _T_5045; // @[Bitwise.scala 48:55:@4421.4]
  wire [1:0] _GEN_718; // @[Bitwise.scala 48:55:@4422.4]
  wire [2:0] _T_5046; // @[Bitwise.scala 48:55:@4422.4]
  wire [2:0] _GEN_719; // @[Bitwise.scala 48:55:@4423.4]
  wire [3:0] _T_5047; // @[Bitwise.scala 48:55:@4423.4]
  wire [3:0] _GEN_720; // @[Bitwise.scala 48:55:@4424.4]
  wire [4:0] _T_5048; // @[Bitwise.scala 48:55:@4424.4]
  wire [1:0] _T_5049; // @[Bitwise.scala 48:55:@4425.4]
  wire [1:0] _T_5050; // @[Bitwise.scala 48:55:@4426.4]
  wire [1:0] _GEN_721; // @[Bitwise.scala 48:55:@4427.4]
  wire [2:0] _T_5051; // @[Bitwise.scala 48:55:@4427.4]
  wire [2:0] _GEN_722; // @[Bitwise.scala 48:55:@4428.4]
  wire [3:0] _T_5052; // @[Bitwise.scala 48:55:@4428.4]
  wire [1:0] _T_5053; // @[Bitwise.scala 48:55:@4429.4]
  wire [1:0] _T_5054; // @[Bitwise.scala 48:55:@4430.4]
  wire [1:0] _GEN_723; // @[Bitwise.scala 48:55:@4431.4]
  wire [2:0] _T_5055; // @[Bitwise.scala 48:55:@4431.4]
  wire [2:0] _GEN_724; // @[Bitwise.scala 48:55:@4432.4]
  wire [3:0] _T_5056; // @[Bitwise.scala 48:55:@4432.4]
  wire [4:0] _T_5057; // @[Bitwise.scala 48:55:@4433.4]
  wire [5:0] _T_5058; // @[Bitwise.scala 48:55:@4434.4]
  wire [1:0] _T_5059; // @[Bitwise.scala 48:55:@4435.4]
  wire [1:0] _T_5060; // @[Bitwise.scala 48:55:@4436.4]
  wire [1:0] _GEN_725; // @[Bitwise.scala 48:55:@4437.4]
  wire [2:0] _T_5061; // @[Bitwise.scala 48:55:@4437.4]
  wire [2:0] _GEN_726; // @[Bitwise.scala 48:55:@4438.4]
  wire [3:0] _T_5062; // @[Bitwise.scala 48:55:@4438.4]
  wire [1:0] _T_5063; // @[Bitwise.scala 48:55:@4439.4]
  wire [1:0] _T_5064; // @[Bitwise.scala 48:55:@4440.4]
  wire [1:0] _GEN_727; // @[Bitwise.scala 48:55:@4441.4]
  wire [2:0] _T_5065; // @[Bitwise.scala 48:55:@4441.4]
  wire [2:0] _GEN_728; // @[Bitwise.scala 48:55:@4442.4]
  wire [3:0] _T_5066; // @[Bitwise.scala 48:55:@4442.4]
  wire [4:0] _T_5067; // @[Bitwise.scala 48:55:@4443.4]
  wire [1:0] _T_5068; // @[Bitwise.scala 48:55:@4444.4]
  wire [1:0] _T_5069; // @[Bitwise.scala 48:55:@4445.4]
  wire [1:0] _GEN_729; // @[Bitwise.scala 48:55:@4446.4]
  wire [2:0] _T_5070; // @[Bitwise.scala 48:55:@4446.4]
  wire [2:0] _GEN_730; // @[Bitwise.scala 48:55:@4447.4]
  wire [3:0] _T_5071; // @[Bitwise.scala 48:55:@4447.4]
  wire [1:0] _T_5072; // @[Bitwise.scala 48:55:@4448.4]
  wire [1:0] _T_5073; // @[Bitwise.scala 48:55:@4449.4]
  wire [1:0] _GEN_731; // @[Bitwise.scala 48:55:@4450.4]
  wire [2:0] _T_5074; // @[Bitwise.scala 48:55:@4450.4]
  wire [2:0] _GEN_732; // @[Bitwise.scala 48:55:@4451.4]
  wire [3:0] _T_5075; // @[Bitwise.scala 48:55:@4451.4]
  wire [4:0] _T_5076; // @[Bitwise.scala 48:55:@4452.4]
  wire [5:0] _T_5077; // @[Bitwise.scala 48:55:@4453.4]
  wire [6:0] _T_5078; // @[Bitwise.scala 48:55:@4454.4]
  wire [39:0] _T_5142; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4519.4]
  wire  _T_5143; // @[Bitwise.scala 50:65:@4520.4]
  wire  _T_5144; // @[Bitwise.scala 50:65:@4521.4]
  wire  _T_5145; // @[Bitwise.scala 50:65:@4522.4]
  wire  _T_5146; // @[Bitwise.scala 50:65:@4523.4]
  wire  _T_5147; // @[Bitwise.scala 50:65:@4524.4]
  wire  _T_5148; // @[Bitwise.scala 50:65:@4525.4]
  wire  _T_5149; // @[Bitwise.scala 50:65:@4526.4]
  wire  _T_5150; // @[Bitwise.scala 50:65:@4527.4]
  wire  _T_5151; // @[Bitwise.scala 50:65:@4528.4]
  wire  _T_5152; // @[Bitwise.scala 50:65:@4529.4]
  wire  _T_5153; // @[Bitwise.scala 50:65:@4530.4]
  wire  _T_5154; // @[Bitwise.scala 50:65:@4531.4]
  wire  _T_5155; // @[Bitwise.scala 50:65:@4532.4]
  wire  _T_5156; // @[Bitwise.scala 50:65:@4533.4]
  wire  _T_5157; // @[Bitwise.scala 50:65:@4534.4]
  wire  _T_5158; // @[Bitwise.scala 50:65:@4535.4]
  wire  _T_5159; // @[Bitwise.scala 50:65:@4536.4]
  wire  _T_5160; // @[Bitwise.scala 50:65:@4537.4]
  wire  _T_5161; // @[Bitwise.scala 50:65:@4538.4]
  wire  _T_5162; // @[Bitwise.scala 50:65:@4539.4]
  wire  _T_5163; // @[Bitwise.scala 50:65:@4540.4]
  wire  _T_5164; // @[Bitwise.scala 50:65:@4541.4]
  wire  _T_5165; // @[Bitwise.scala 50:65:@4542.4]
  wire  _T_5166; // @[Bitwise.scala 50:65:@4543.4]
  wire  _T_5167; // @[Bitwise.scala 50:65:@4544.4]
  wire  _T_5168; // @[Bitwise.scala 50:65:@4545.4]
  wire  _T_5169; // @[Bitwise.scala 50:65:@4546.4]
  wire  _T_5170; // @[Bitwise.scala 50:65:@4547.4]
  wire  _T_5171; // @[Bitwise.scala 50:65:@4548.4]
  wire  _T_5172; // @[Bitwise.scala 50:65:@4549.4]
  wire  _T_5173; // @[Bitwise.scala 50:65:@4550.4]
  wire  _T_5174; // @[Bitwise.scala 50:65:@4551.4]
  wire  _T_5175; // @[Bitwise.scala 50:65:@4552.4]
  wire  _T_5176; // @[Bitwise.scala 50:65:@4553.4]
  wire  _T_5177; // @[Bitwise.scala 50:65:@4554.4]
  wire  _T_5178; // @[Bitwise.scala 50:65:@4555.4]
  wire  _T_5179; // @[Bitwise.scala 50:65:@4556.4]
  wire  _T_5180; // @[Bitwise.scala 50:65:@4557.4]
  wire  _T_5181; // @[Bitwise.scala 50:65:@4558.4]
  wire  _T_5182; // @[Bitwise.scala 50:65:@4559.4]
  wire [1:0] _T_5183; // @[Bitwise.scala 48:55:@4560.4]
  wire [1:0] _T_5184; // @[Bitwise.scala 48:55:@4561.4]
  wire [1:0] _GEN_733; // @[Bitwise.scala 48:55:@4562.4]
  wire [2:0] _T_5185; // @[Bitwise.scala 48:55:@4562.4]
  wire [2:0] _GEN_734; // @[Bitwise.scala 48:55:@4563.4]
  wire [3:0] _T_5186; // @[Bitwise.scala 48:55:@4563.4]
  wire [1:0] _T_5187; // @[Bitwise.scala 48:55:@4564.4]
  wire [1:0] _T_5188; // @[Bitwise.scala 48:55:@4565.4]
  wire [1:0] _GEN_735; // @[Bitwise.scala 48:55:@4566.4]
  wire [2:0] _T_5189; // @[Bitwise.scala 48:55:@4566.4]
  wire [2:0] _GEN_736; // @[Bitwise.scala 48:55:@4567.4]
  wire [3:0] _T_5190; // @[Bitwise.scala 48:55:@4567.4]
  wire [4:0] _T_5191; // @[Bitwise.scala 48:55:@4568.4]
  wire [1:0] _T_5192; // @[Bitwise.scala 48:55:@4569.4]
  wire [1:0] _T_5193; // @[Bitwise.scala 48:55:@4570.4]
  wire [1:0] _GEN_737; // @[Bitwise.scala 48:55:@4571.4]
  wire [2:0] _T_5194; // @[Bitwise.scala 48:55:@4571.4]
  wire [2:0] _GEN_738; // @[Bitwise.scala 48:55:@4572.4]
  wire [3:0] _T_5195; // @[Bitwise.scala 48:55:@4572.4]
  wire [1:0] _T_5196; // @[Bitwise.scala 48:55:@4573.4]
  wire [1:0] _T_5197; // @[Bitwise.scala 48:55:@4574.4]
  wire [1:0] _GEN_739; // @[Bitwise.scala 48:55:@4575.4]
  wire [2:0] _T_5198; // @[Bitwise.scala 48:55:@4575.4]
  wire [2:0] _GEN_740; // @[Bitwise.scala 48:55:@4576.4]
  wire [3:0] _T_5199; // @[Bitwise.scala 48:55:@4576.4]
  wire [4:0] _T_5200; // @[Bitwise.scala 48:55:@4577.4]
  wire [5:0] _T_5201; // @[Bitwise.scala 48:55:@4578.4]
  wire [1:0] _T_5202; // @[Bitwise.scala 48:55:@4579.4]
  wire [1:0] _T_5203; // @[Bitwise.scala 48:55:@4580.4]
  wire [1:0] _GEN_741; // @[Bitwise.scala 48:55:@4581.4]
  wire [2:0] _T_5204; // @[Bitwise.scala 48:55:@4581.4]
  wire [2:0] _GEN_742; // @[Bitwise.scala 48:55:@4582.4]
  wire [3:0] _T_5205; // @[Bitwise.scala 48:55:@4582.4]
  wire [1:0] _T_5206; // @[Bitwise.scala 48:55:@4583.4]
  wire [1:0] _T_5207; // @[Bitwise.scala 48:55:@4584.4]
  wire [1:0] _GEN_743; // @[Bitwise.scala 48:55:@4585.4]
  wire [2:0] _T_5208; // @[Bitwise.scala 48:55:@4585.4]
  wire [2:0] _GEN_744; // @[Bitwise.scala 48:55:@4586.4]
  wire [3:0] _T_5209; // @[Bitwise.scala 48:55:@4586.4]
  wire [4:0] _T_5210; // @[Bitwise.scala 48:55:@4587.4]
  wire [1:0] _T_5211; // @[Bitwise.scala 48:55:@4588.4]
  wire [1:0] _T_5212; // @[Bitwise.scala 48:55:@4589.4]
  wire [1:0] _GEN_745; // @[Bitwise.scala 48:55:@4590.4]
  wire [2:0] _T_5213; // @[Bitwise.scala 48:55:@4590.4]
  wire [2:0] _GEN_746; // @[Bitwise.scala 48:55:@4591.4]
  wire [3:0] _T_5214; // @[Bitwise.scala 48:55:@4591.4]
  wire [1:0] _T_5215; // @[Bitwise.scala 48:55:@4592.4]
  wire [1:0] _T_5216; // @[Bitwise.scala 48:55:@4593.4]
  wire [1:0] _GEN_747; // @[Bitwise.scala 48:55:@4594.4]
  wire [2:0] _T_5217; // @[Bitwise.scala 48:55:@4594.4]
  wire [2:0] _GEN_748; // @[Bitwise.scala 48:55:@4595.4]
  wire [3:0] _T_5218; // @[Bitwise.scala 48:55:@4595.4]
  wire [4:0] _T_5219; // @[Bitwise.scala 48:55:@4596.4]
  wire [5:0] _T_5220; // @[Bitwise.scala 48:55:@4597.4]
  wire [6:0] _T_5221; // @[Bitwise.scala 48:55:@4598.4]
  wire [40:0] _T_5285; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4663.4]
  wire  _T_5286; // @[Bitwise.scala 50:65:@4664.4]
  wire  _T_5287; // @[Bitwise.scala 50:65:@4665.4]
  wire  _T_5288; // @[Bitwise.scala 50:65:@4666.4]
  wire  _T_5289; // @[Bitwise.scala 50:65:@4667.4]
  wire  _T_5290; // @[Bitwise.scala 50:65:@4668.4]
  wire  _T_5291; // @[Bitwise.scala 50:65:@4669.4]
  wire  _T_5292; // @[Bitwise.scala 50:65:@4670.4]
  wire  _T_5293; // @[Bitwise.scala 50:65:@4671.4]
  wire  _T_5294; // @[Bitwise.scala 50:65:@4672.4]
  wire  _T_5295; // @[Bitwise.scala 50:65:@4673.4]
  wire  _T_5296; // @[Bitwise.scala 50:65:@4674.4]
  wire  _T_5297; // @[Bitwise.scala 50:65:@4675.4]
  wire  _T_5298; // @[Bitwise.scala 50:65:@4676.4]
  wire  _T_5299; // @[Bitwise.scala 50:65:@4677.4]
  wire  _T_5300; // @[Bitwise.scala 50:65:@4678.4]
  wire  _T_5301; // @[Bitwise.scala 50:65:@4679.4]
  wire  _T_5302; // @[Bitwise.scala 50:65:@4680.4]
  wire  _T_5303; // @[Bitwise.scala 50:65:@4681.4]
  wire  _T_5304; // @[Bitwise.scala 50:65:@4682.4]
  wire  _T_5305; // @[Bitwise.scala 50:65:@4683.4]
  wire  _T_5306; // @[Bitwise.scala 50:65:@4684.4]
  wire  _T_5307; // @[Bitwise.scala 50:65:@4685.4]
  wire  _T_5308; // @[Bitwise.scala 50:65:@4686.4]
  wire  _T_5309; // @[Bitwise.scala 50:65:@4687.4]
  wire  _T_5310; // @[Bitwise.scala 50:65:@4688.4]
  wire  _T_5311; // @[Bitwise.scala 50:65:@4689.4]
  wire  _T_5312; // @[Bitwise.scala 50:65:@4690.4]
  wire  _T_5313; // @[Bitwise.scala 50:65:@4691.4]
  wire  _T_5314; // @[Bitwise.scala 50:65:@4692.4]
  wire  _T_5315; // @[Bitwise.scala 50:65:@4693.4]
  wire  _T_5316; // @[Bitwise.scala 50:65:@4694.4]
  wire  _T_5317; // @[Bitwise.scala 50:65:@4695.4]
  wire  _T_5318; // @[Bitwise.scala 50:65:@4696.4]
  wire  _T_5319; // @[Bitwise.scala 50:65:@4697.4]
  wire  _T_5320; // @[Bitwise.scala 50:65:@4698.4]
  wire  _T_5321; // @[Bitwise.scala 50:65:@4699.4]
  wire  _T_5322; // @[Bitwise.scala 50:65:@4700.4]
  wire  _T_5323; // @[Bitwise.scala 50:65:@4701.4]
  wire  _T_5324; // @[Bitwise.scala 50:65:@4702.4]
  wire  _T_5325; // @[Bitwise.scala 50:65:@4703.4]
  wire  _T_5326; // @[Bitwise.scala 50:65:@4704.4]
  wire [1:0] _T_5327; // @[Bitwise.scala 48:55:@4705.4]
  wire [1:0] _T_5328; // @[Bitwise.scala 48:55:@4706.4]
  wire [1:0] _GEN_749; // @[Bitwise.scala 48:55:@4707.4]
  wire [2:0] _T_5329; // @[Bitwise.scala 48:55:@4707.4]
  wire [2:0] _GEN_750; // @[Bitwise.scala 48:55:@4708.4]
  wire [3:0] _T_5330; // @[Bitwise.scala 48:55:@4708.4]
  wire [1:0] _T_5331; // @[Bitwise.scala 48:55:@4709.4]
  wire [1:0] _T_5332; // @[Bitwise.scala 48:55:@4710.4]
  wire [1:0] _GEN_751; // @[Bitwise.scala 48:55:@4711.4]
  wire [2:0] _T_5333; // @[Bitwise.scala 48:55:@4711.4]
  wire [2:0] _GEN_752; // @[Bitwise.scala 48:55:@4712.4]
  wire [3:0] _T_5334; // @[Bitwise.scala 48:55:@4712.4]
  wire [4:0] _T_5335; // @[Bitwise.scala 48:55:@4713.4]
  wire [1:0] _T_5336; // @[Bitwise.scala 48:55:@4714.4]
  wire [1:0] _T_5337; // @[Bitwise.scala 48:55:@4715.4]
  wire [1:0] _GEN_753; // @[Bitwise.scala 48:55:@4716.4]
  wire [2:0] _T_5338; // @[Bitwise.scala 48:55:@4716.4]
  wire [2:0] _GEN_754; // @[Bitwise.scala 48:55:@4717.4]
  wire [3:0] _T_5339; // @[Bitwise.scala 48:55:@4717.4]
  wire [1:0] _T_5340; // @[Bitwise.scala 48:55:@4718.4]
  wire [1:0] _T_5341; // @[Bitwise.scala 48:55:@4719.4]
  wire [1:0] _GEN_755; // @[Bitwise.scala 48:55:@4720.4]
  wire [2:0] _T_5342; // @[Bitwise.scala 48:55:@4720.4]
  wire [2:0] _GEN_756; // @[Bitwise.scala 48:55:@4721.4]
  wire [3:0] _T_5343; // @[Bitwise.scala 48:55:@4721.4]
  wire [4:0] _T_5344; // @[Bitwise.scala 48:55:@4722.4]
  wire [5:0] _T_5345; // @[Bitwise.scala 48:55:@4723.4]
  wire [1:0] _T_5346; // @[Bitwise.scala 48:55:@4724.4]
  wire [1:0] _T_5347; // @[Bitwise.scala 48:55:@4725.4]
  wire [1:0] _GEN_757; // @[Bitwise.scala 48:55:@4726.4]
  wire [2:0] _T_5348; // @[Bitwise.scala 48:55:@4726.4]
  wire [2:0] _GEN_758; // @[Bitwise.scala 48:55:@4727.4]
  wire [3:0] _T_5349; // @[Bitwise.scala 48:55:@4727.4]
  wire [1:0] _T_5350; // @[Bitwise.scala 48:55:@4728.4]
  wire [1:0] _T_5351; // @[Bitwise.scala 48:55:@4729.4]
  wire [1:0] _GEN_759; // @[Bitwise.scala 48:55:@4730.4]
  wire [2:0] _T_5352; // @[Bitwise.scala 48:55:@4730.4]
  wire [2:0] _GEN_760; // @[Bitwise.scala 48:55:@4731.4]
  wire [3:0] _T_5353; // @[Bitwise.scala 48:55:@4731.4]
  wire [4:0] _T_5354; // @[Bitwise.scala 48:55:@4732.4]
  wire [1:0] _T_5355; // @[Bitwise.scala 48:55:@4733.4]
  wire [1:0] _T_5356; // @[Bitwise.scala 48:55:@4734.4]
  wire [1:0] _GEN_761; // @[Bitwise.scala 48:55:@4735.4]
  wire [2:0] _T_5357; // @[Bitwise.scala 48:55:@4735.4]
  wire [2:0] _GEN_762; // @[Bitwise.scala 48:55:@4736.4]
  wire [3:0] _T_5358; // @[Bitwise.scala 48:55:@4736.4]
  wire [1:0] _T_5359; // @[Bitwise.scala 48:55:@4737.4]
  wire [1:0] _GEN_763; // @[Bitwise.scala 48:55:@4738.4]
  wire [2:0] _T_5360; // @[Bitwise.scala 48:55:@4738.4]
  wire [1:0] _T_5361; // @[Bitwise.scala 48:55:@4739.4]
  wire [1:0] _GEN_764; // @[Bitwise.scala 48:55:@4740.4]
  wire [2:0] _T_5362; // @[Bitwise.scala 48:55:@4740.4]
  wire [3:0] _T_5363; // @[Bitwise.scala 48:55:@4741.4]
  wire [4:0] _T_5364; // @[Bitwise.scala 48:55:@4742.4]
  wire [5:0] _T_5365; // @[Bitwise.scala 48:55:@4743.4]
  wire [6:0] _T_5366; // @[Bitwise.scala 48:55:@4744.4]
  wire [41:0] _T_5430; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4809.4]
  wire  _T_5431; // @[Bitwise.scala 50:65:@4810.4]
  wire  _T_5432; // @[Bitwise.scala 50:65:@4811.4]
  wire  _T_5433; // @[Bitwise.scala 50:65:@4812.4]
  wire  _T_5434; // @[Bitwise.scala 50:65:@4813.4]
  wire  _T_5435; // @[Bitwise.scala 50:65:@4814.4]
  wire  _T_5436; // @[Bitwise.scala 50:65:@4815.4]
  wire  _T_5437; // @[Bitwise.scala 50:65:@4816.4]
  wire  _T_5438; // @[Bitwise.scala 50:65:@4817.4]
  wire  _T_5439; // @[Bitwise.scala 50:65:@4818.4]
  wire  _T_5440; // @[Bitwise.scala 50:65:@4819.4]
  wire  _T_5441; // @[Bitwise.scala 50:65:@4820.4]
  wire  _T_5442; // @[Bitwise.scala 50:65:@4821.4]
  wire  _T_5443; // @[Bitwise.scala 50:65:@4822.4]
  wire  _T_5444; // @[Bitwise.scala 50:65:@4823.4]
  wire  _T_5445; // @[Bitwise.scala 50:65:@4824.4]
  wire  _T_5446; // @[Bitwise.scala 50:65:@4825.4]
  wire  _T_5447; // @[Bitwise.scala 50:65:@4826.4]
  wire  _T_5448; // @[Bitwise.scala 50:65:@4827.4]
  wire  _T_5449; // @[Bitwise.scala 50:65:@4828.4]
  wire  _T_5450; // @[Bitwise.scala 50:65:@4829.4]
  wire  _T_5451; // @[Bitwise.scala 50:65:@4830.4]
  wire  _T_5452; // @[Bitwise.scala 50:65:@4831.4]
  wire  _T_5453; // @[Bitwise.scala 50:65:@4832.4]
  wire  _T_5454; // @[Bitwise.scala 50:65:@4833.4]
  wire  _T_5455; // @[Bitwise.scala 50:65:@4834.4]
  wire  _T_5456; // @[Bitwise.scala 50:65:@4835.4]
  wire  _T_5457; // @[Bitwise.scala 50:65:@4836.4]
  wire  _T_5458; // @[Bitwise.scala 50:65:@4837.4]
  wire  _T_5459; // @[Bitwise.scala 50:65:@4838.4]
  wire  _T_5460; // @[Bitwise.scala 50:65:@4839.4]
  wire  _T_5461; // @[Bitwise.scala 50:65:@4840.4]
  wire  _T_5462; // @[Bitwise.scala 50:65:@4841.4]
  wire  _T_5463; // @[Bitwise.scala 50:65:@4842.4]
  wire  _T_5464; // @[Bitwise.scala 50:65:@4843.4]
  wire  _T_5465; // @[Bitwise.scala 50:65:@4844.4]
  wire  _T_5466; // @[Bitwise.scala 50:65:@4845.4]
  wire  _T_5467; // @[Bitwise.scala 50:65:@4846.4]
  wire  _T_5468; // @[Bitwise.scala 50:65:@4847.4]
  wire  _T_5469; // @[Bitwise.scala 50:65:@4848.4]
  wire  _T_5470; // @[Bitwise.scala 50:65:@4849.4]
  wire  _T_5471; // @[Bitwise.scala 50:65:@4850.4]
  wire  _T_5472; // @[Bitwise.scala 50:65:@4851.4]
  wire [1:0] _T_5473; // @[Bitwise.scala 48:55:@4852.4]
  wire [1:0] _T_5474; // @[Bitwise.scala 48:55:@4853.4]
  wire [1:0] _GEN_765; // @[Bitwise.scala 48:55:@4854.4]
  wire [2:0] _T_5475; // @[Bitwise.scala 48:55:@4854.4]
  wire [2:0] _GEN_766; // @[Bitwise.scala 48:55:@4855.4]
  wire [3:0] _T_5476; // @[Bitwise.scala 48:55:@4855.4]
  wire [1:0] _T_5477; // @[Bitwise.scala 48:55:@4856.4]
  wire [1:0] _T_5478; // @[Bitwise.scala 48:55:@4857.4]
  wire [1:0] _GEN_767; // @[Bitwise.scala 48:55:@4858.4]
  wire [2:0] _T_5479; // @[Bitwise.scala 48:55:@4858.4]
  wire [2:0] _GEN_768; // @[Bitwise.scala 48:55:@4859.4]
  wire [3:0] _T_5480; // @[Bitwise.scala 48:55:@4859.4]
  wire [4:0] _T_5481; // @[Bitwise.scala 48:55:@4860.4]
  wire [1:0] _T_5482; // @[Bitwise.scala 48:55:@4861.4]
  wire [1:0] _T_5483; // @[Bitwise.scala 48:55:@4862.4]
  wire [1:0] _GEN_769; // @[Bitwise.scala 48:55:@4863.4]
  wire [2:0] _T_5484; // @[Bitwise.scala 48:55:@4863.4]
  wire [2:0] _GEN_770; // @[Bitwise.scala 48:55:@4864.4]
  wire [3:0] _T_5485; // @[Bitwise.scala 48:55:@4864.4]
  wire [1:0] _T_5486; // @[Bitwise.scala 48:55:@4865.4]
  wire [1:0] _GEN_771; // @[Bitwise.scala 48:55:@4866.4]
  wire [2:0] _T_5487; // @[Bitwise.scala 48:55:@4866.4]
  wire [1:0] _T_5488; // @[Bitwise.scala 48:55:@4867.4]
  wire [1:0] _GEN_772; // @[Bitwise.scala 48:55:@4868.4]
  wire [2:0] _T_5489; // @[Bitwise.scala 48:55:@4868.4]
  wire [3:0] _T_5490; // @[Bitwise.scala 48:55:@4869.4]
  wire [4:0] _T_5491; // @[Bitwise.scala 48:55:@4870.4]
  wire [5:0] _T_5492; // @[Bitwise.scala 48:55:@4871.4]
  wire [1:0] _T_5493; // @[Bitwise.scala 48:55:@4872.4]
  wire [1:0] _T_5494; // @[Bitwise.scala 48:55:@4873.4]
  wire [1:0] _GEN_773; // @[Bitwise.scala 48:55:@4874.4]
  wire [2:0] _T_5495; // @[Bitwise.scala 48:55:@4874.4]
  wire [2:0] _GEN_774; // @[Bitwise.scala 48:55:@4875.4]
  wire [3:0] _T_5496; // @[Bitwise.scala 48:55:@4875.4]
  wire [1:0] _T_5497; // @[Bitwise.scala 48:55:@4876.4]
  wire [1:0] _T_5498; // @[Bitwise.scala 48:55:@4877.4]
  wire [1:0] _GEN_775; // @[Bitwise.scala 48:55:@4878.4]
  wire [2:0] _T_5499; // @[Bitwise.scala 48:55:@4878.4]
  wire [2:0] _GEN_776; // @[Bitwise.scala 48:55:@4879.4]
  wire [3:0] _T_5500; // @[Bitwise.scala 48:55:@4879.4]
  wire [4:0] _T_5501; // @[Bitwise.scala 48:55:@4880.4]
  wire [1:0] _T_5502; // @[Bitwise.scala 48:55:@4881.4]
  wire [1:0] _T_5503; // @[Bitwise.scala 48:55:@4882.4]
  wire [1:0] _GEN_777; // @[Bitwise.scala 48:55:@4883.4]
  wire [2:0] _T_5504; // @[Bitwise.scala 48:55:@4883.4]
  wire [2:0] _GEN_778; // @[Bitwise.scala 48:55:@4884.4]
  wire [3:0] _T_5505; // @[Bitwise.scala 48:55:@4884.4]
  wire [1:0] _T_5506; // @[Bitwise.scala 48:55:@4885.4]
  wire [1:0] _GEN_779; // @[Bitwise.scala 48:55:@4886.4]
  wire [2:0] _T_5507; // @[Bitwise.scala 48:55:@4886.4]
  wire [1:0] _T_5508; // @[Bitwise.scala 48:55:@4887.4]
  wire [1:0] _GEN_780; // @[Bitwise.scala 48:55:@4888.4]
  wire [2:0] _T_5509; // @[Bitwise.scala 48:55:@4888.4]
  wire [3:0] _T_5510; // @[Bitwise.scala 48:55:@4889.4]
  wire [4:0] _T_5511; // @[Bitwise.scala 48:55:@4890.4]
  wire [5:0] _T_5512; // @[Bitwise.scala 48:55:@4891.4]
  wire [6:0] _T_5513; // @[Bitwise.scala 48:55:@4892.4]
  wire [42:0] _T_5577; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4957.4]
  wire  _T_5578; // @[Bitwise.scala 50:65:@4958.4]
  wire  _T_5579; // @[Bitwise.scala 50:65:@4959.4]
  wire  _T_5580; // @[Bitwise.scala 50:65:@4960.4]
  wire  _T_5581; // @[Bitwise.scala 50:65:@4961.4]
  wire  _T_5582; // @[Bitwise.scala 50:65:@4962.4]
  wire  _T_5583; // @[Bitwise.scala 50:65:@4963.4]
  wire  _T_5584; // @[Bitwise.scala 50:65:@4964.4]
  wire  _T_5585; // @[Bitwise.scala 50:65:@4965.4]
  wire  _T_5586; // @[Bitwise.scala 50:65:@4966.4]
  wire  _T_5587; // @[Bitwise.scala 50:65:@4967.4]
  wire  _T_5588; // @[Bitwise.scala 50:65:@4968.4]
  wire  _T_5589; // @[Bitwise.scala 50:65:@4969.4]
  wire  _T_5590; // @[Bitwise.scala 50:65:@4970.4]
  wire  _T_5591; // @[Bitwise.scala 50:65:@4971.4]
  wire  _T_5592; // @[Bitwise.scala 50:65:@4972.4]
  wire  _T_5593; // @[Bitwise.scala 50:65:@4973.4]
  wire  _T_5594; // @[Bitwise.scala 50:65:@4974.4]
  wire  _T_5595; // @[Bitwise.scala 50:65:@4975.4]
  wire  _T_5596; // @[Bitwise.scala 50:65:@4976.4]
  wire  _T_5597; // @[Bitwise.scala 50:65:@4977.4]
  wire  _T_5598; // @[Bitwise.scala 50:65:@4978.4]
  wire  _T_5599; // @[Bitwise.scala 50:65:@4979.4]
  wire  _T_5600; // @[Bitwise.scala 50:65:@4980.4]
  wire  _T_5601; // @[Bitwise.scala 50:65:@4981.4]
  wire  _T_5602; // @[Bitwise.scala 50:65:@4982.4]
  wire  _T_5603; // @[Bitwise.scala 50:65:@4983.4]
  wire  _T_5604; // @[Bitwise.scala 50:65:@4984.4]
  wire  _T_5605; // @[Bitwise.scala 50:65:@4985.4]
  wire  _T_5606; // @[Bitwise.scala 50:65:@4986.4]
  wire  _T_5607; // @[Bitwise.scala 50:65:@4987.4]
  wire  _T_5608; // @[Bitwise.scala 50:65:@4988.4]
  wire  _T_5609; // @[Bitwise.scala 50:65:@4989.4]
  wire  _T_5610; // @[Bitwise.scala 50:65:@4990.4]
  wire  _T_5611; // @[Bitwise.scala 50:65:@4991.4]
  wire  _T_5612; // @[Bitwise.scala 50:65:@4992.4]
  wire  _T_5613; // @[Bitwise.scala 50:65:@4993.4]
  wire  _T_5614; // @[Bitwise.scala 50:65:@4994.4]
  wire  _T_5615; // @[Bitwise.scala 50:65:@4995.4]
  wire  _T_5616; // @[Bitwise.scala 50:65:@4996.4]
  wire  _T_5617; // @[Bitwise.scala 50:65:@4997.4]
  wire  _T_5618; // @[Bitwise.scala 50:65:@4998.4]
  wire  _T_5619; // @[Bitwise.scala 50:65:@4999.4]
  wire  _T_5620; // @[Bitwise.scala 50:65:@5000.4]
  wire [1:0] _T_5621; // @[Bitwise.scala 48:55:@5001.4]
  wire [1:0] _T_5622; // @[Bitwise.scala 48:55:@5002.4]
  wire [1:0] _GEN_781; // @[Bitwise.scala 48:55:@5003.4]
  wire [2:0] _T_5623; // @[Bitwise.scala 48:55:@5003.4]
  wire [2:0] _GEN_782; // @[Bitwise.scala 48:55:@5004.4]
  wire [3:0] _T_5624; // @[Bitwise.scala 48:55:@5004.4]
  wire [1:0] _T_5625; // @[Bitwise.scala 48:55:@5005.4]
  wire [1:0] _T_5626; // @[Bitwise.scala 48:55:@5006.4]
  wire [1:0] _GEN_783; // @[Bitwise.scala 48:55:@5007.4]
  wire [2:0] _T_5627; // @[Bitwise.scala 48:55:@5007.4]
  wire [2:0] _GEN_784; // @[Bitwise.scala 48:55:@5008.4]
  wire [3:0] _T_5628; // @[Bitwise.scala 48:55:@5008.4]
  wire [4:0] _T_5629; // @[Bitwise.scala 48:55:@5009.4]
  wire [1:0] _T_5630; // @[Bitwise.scala 48:55:@5010.4]
  wire [1:0] _T_5631; // @[Bitwise.scala 48:55:@5011.4]
  wire [1:0] _GEN_785; // @[Bitwise.scala 48:55:@5012.4]
  wire [2:0] _T_5632; // @[Bitwise.scala 48:55:@5012.4]
  wire [2:0] _GEN_786; // @[Bitwise.scala 48:55:@5013.4]
  wire [3:0] _T_5633; // @[Bitwise.scala 48:55:@5013.4]
  wire [1:0] _T_5634; // @[Bitwise.scala 48:55:@5014.4]
  wire [1:0] _GEN_787; // @[Bitwise.scala 48:55:@5015.4]
  wire [2:0] _T_5635; // @[Bitwise.scala 48:55:@5015.4]
  wire [1:0] _T_5636; // @[Bitwise.scala 48:55:@5016.4]
  wire [1:0] _GEN_788; // @[Bitwise.scala 48:55:@5017.4]
  wire [2:0] _T_5637; // @[Bitwise.scala 48:55:@5017.4]
  wire [3:0] _T_5638; // @[Bitwise.scala 48:55:@5018.4]
  wire [4:0] _T_5639; // @[Bitwise.scala 48:55:@5019.4]
  wire [5:0] _T_5640; // @[Bitwise.scala 48:55:@5020.4]
  wire [1:0] _T_5641; // @[Bitwise.scala 48:55:@5021.4]
  wire [1:0] _T_5642; // @[Bitwise.scala 48:55:@5022.4]
  wire [1:0] _GEN_789; // @[Bitwise.scala 48:55:@5023.4]
  wire [2:0] _T_5643; // @[Bitwise.scala 48:55:@5023.4]
  wire [2:0] _GEN_790; // @[Bitwise.scala 48:55:@5024.4]
  wire [3:0] _T_5644; // @[Bitwise.scala 48:55:@5024.4]
  wire [1:0] _T_5645; // @[Bitwise.scala 48:55:@5025.4]
  wire [1:0] _GEN_791; // @[Bitwise.scala 48:55:@5026.4]
  wire [2:0] _T_5646; // @[Bitwise.scala 48:55:@5026.4]
  wire [1:0] _T_5647; // @[Bitwise.scala 48:55:@5027.4]
  wire [1:0] _GEN_792; // @[Bitwise.scala 48:55:@5028.4]
  wire [2:0] _T_5648; // @[Bitwise.scala 48:55:@5028.4]
  wire [3:0] _T_5649; // @[Bitwise.scala 48:55:@5029.4]
  wire [4:0] _T_5650; // @[Bitwise.scala 48:55:@5030.4]
  wire [1:0] _T_5651; // @[Bitwise.scala 48:55:@5031.4]
  wire [1:0] _T_5652; // @[Bitwise.scala 48:55:@5032.4]
  wire [1:0] _GEN_793; // @[Bitwise.scala 48:55:@5033.4]
  wire [2:0] _T_5653; // @[Bitwise.scala 48:55:@5033.4]
  wire [2:0] _GEN_794; // @[Bitwise.scala 48:55:@5034.4]
  wire [3:0] _T_5654; // @[Bitwise.scala 48:55:@5034.4]
  wire [1:0] _T_5655; // @[Bitwise.scala 48:55:@5035.4]
  wire [1:0] _GEN_795; // @[Bitwise.scala 48:55:@5036.4]
  wire [2:0] _T_5656; // @[Bitwise.scala 48:55:@5036.4]
  wire [1:0] _T_5657; // @[Bitwise.scala 48:55:@5037.4]
  wire [1:0] _GEN_796; // @[Bitwise.scala 48:55:@5038.4]
  wire [2:0] _T_5658; // @[Bitwise.scala 48:55:@5038.4]
  wire [3:0] _T_5659; // @[Bitwise.scala 48:55:@5039.4]
  wire [4:0] _T_5660; // @[Bitwise.scala 48:55:@5040.4]
  wire [5:0] _T_5661; // @[Bitwise.scala 48:55:@5041.4]
  wire [6:0] _T_5662; // @[Bitwise.scala 48:55:@5042.4]
  wire [43:0] _T_5726; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5107.4]
  wire  _T_5727; // @[Bitwise.scala 50:65:@5108.4]
  wire  _T_5728; // @[Bitwise.scala 50:65:@5109.4]
  wire  _T_5729; // @[Bitwise.scala 50:65:@5110.4]
  wire  _T_5730; // @[Bitwise.scala 50:65:@5111.4]
  wire  _T_5731; // @[Bitwise.scala 50:65:@5112.4]
  wire  _T_5732; // @[Bitwise.scala 50:65:@5113.4]
  wire  _T_5733; // @[Bitwise.scala 50:65:@5114.4]
  wire  _T_5734; // @[Bitwise.scala 50:65:@5115.4]
  wire  _T_5735; // @[Bitwise.scala 50:65:@5116.4]
  wire  _T_5736; // @[Bitwise.scala 50:65:@5117.4]
  wire  _T_5737; // @[Bitwise.scala 50:65:@5118.4]
  wire  _T_5738; // @[Bitwise.scala 50:65:@5119.4]
  wire  _T_5739; // @[Bitwise.scala 50:65:@5120.4]
  wire  _T_5740; // @[Bitwise.scala 50:65:@5121.4]
  wire  _T_5741; // @[Bitwise.scala 50:65:@5122.4]
  wire  _T_5742; // @[Bitwise.scala 50:65:@5123.4]
  wire  _T_5743; // @[Bitwise.scala 50:65:@5124.4]
  wire  _T_5744; // @[Bitwise.scala 50:65:@5125.4]
  wire  _T_5745; // @[Bitwise.scala 50:65:@5126.4]
  wire  _T_5746; // @[Bitwise.scala 50:65:@5127.4]
  wire  _T_5747; // @[Bitwise.scala 50:65:@5128.4]
  wire  _T_5748; // @[Bitwise.scala 50:65:@5129.4]
  wire  _T_5749; // @[Bitwise.scala 50:65:@5130.4]
  wire  _T_5750; // @[Bitwise.scala 50:65:@5131.4]
  wire  _T_5751; // @[Bitwise.scala 50:65:@5132.4]
  wire  _T_5752; // @[Bitwise.scala 50:65:@5133.4]
  wire  _T_5753; // @[Bitwise.scala 50:65:@5134.4]
  wire  _T_5754; // @[Bitwise.scala 50:65:@5135.4]
  wire  _T_5755; // @[Bitwise.scala 50:65:@5136.4]
  wire  _T_5756; // @[Bitwise.scala 50:65:@5137.4]
  wire  _T_5757; // @[Bitwise.scala 50:65:@5138.4]
  wire  _T_5758; // @[Bitwise.scala 50:65:@5139.4]
  wire  _T_5759; // @[Bitwise.scala 50:65:@5140.4]
  wire  _T_5760; // @[Bitwise.scala 50:65:@5141.4]
  wire  _T_5761; // @[Bitwise.scala 50:65:@5142.4]
  wire  _T_5762; // @[Bitwise.scala 50:65:@5143.4]
  wire  _T_5763; // @[Bitwise.scala 50:65:@5144.4]
  wire  _T_5764; // @[Bitwise.scala 50:65:@5145.4]
  wire  _T_5765; // @[Bitwise.scala 50:65:@5146.4]
  wire  _T_5766; // @[Bitwise.scala 50:65:@5147.4]
  wire  _T_5767; // @[Bitwise.scala 50:65:@5148.4]
  wire  _T_5768; // @[Bitwise.scala 50:65:@5149.4]
  wire  _T_5769; // @[Bitwise.scala 50:65:@5150.4]
  wire  _T_5770; // @[Bitwise.scala 50:65:@5151.4]
  wire [1:0] _T_5771; // @[Bitwise.scala 48:55:@5152.4]
  wire [1:0] _T_5772; // @[Bitwise.scala 48:55:@5153.4]
  wire [1:0] _GEN_797; // @[Bitwise.scala 48:55:@5154.4]
  wire [2:0] _T_5773; // @[Bitwise.scala 48:55:@5154.4]
  wire [2:0] _GEN_798; // @[Bitwise.scala 48:55:@5155.4]
  wire [3:0] _T_5774; // @[Bitwise.scala 48:55:@5155.4]
  wire [1:0] _T_5775; // @[Bitwise.scala 48:55:@5156.4]
  wire [1:0] _GEN_799; // @[Bitwise.scala 48:55:@5157.4]
  wire [2:0] _T_5776; // @[Bitwise.scala 48:55:@5157.4]
  wire [1:0] _T_5777; // @[Bitwise.scala 48:55:@5158.4]
  wire [1:0] _GEN_800; // @[Bitwise.scala 48:55:@5159.4]
  wire [2:0] _T_5778; // @[Bitwise.scala 48:55:@5159.4]
  wire [3:0] _T_5779; // @[Bitwise.scala 48:55:@5160.4]
  wire [4:0] _T_5780; // @[Bitwise.scala 48:55:@5161.4]
  wire [1:0] _T_5781; // @[Bitwise.scala 48:55:@5162.4]
  wire [1:0] _T_5782; // @[Bitwise.scala 48:55:@5163.4]
  wire [1:0] _GEN_801; // @[Bitwise.scala 48:55:@5164.4]
  wire [2:0] _T_5783; // @[Bitwise.scala 48:55:@5164.4]
  wire [2:0] _GEN_802; // @[Bitwise.scala 48:55:@5165.4]
  wire [3:0] _T_5784; // @[Bitwise.scala 48:55:@5165.4]
  wire [1:0] _T_5785; // @[Bitwise.scala 48:55:@5166.4]
  wire [1:0] _GEN_803; // @[Bitwise.scala 48:55:@5167.4]
  wire [2:0] _T_5786; // @[Bitwise.scala 48:55:@5167.4]
  wire [1:0] _T_5787; // @[Bitwise.scala 48:55:@5168.4]
  wire [1:0] _GEN_804; // @[Bitwise.scala 48:55:@5169.4]
  wire [2:0] _T_5788; // @[Bitwise.scala 48:55:@5169.4]
  wire [3:0] _T_5789; // @[Bitwise.scala 48:55:@5170.4]
  wire [4:0] _T_5790; // @[Bitwise.scala 48:55:@5171.4]
  wire [5:0] _T_5791; // @[Bitwise.scala 48:55:@5172.4]
  wire [1:0] _T_5792; // @[Bitwise.scala 48:55:@5173.4]
  wire [1:0] _T_5793; // @[Bitwise.scala 48:55:@5174.4]
  wire [1:0] _GEN_805; // @[Bitwise.scala 48:55:@5175.4]
  wire [2:0] _T_5794; // @[Bitwise.scala 48:55:@5175.4]
  wire [2:0] _GEN_806; // @[Bitwise.scala 48:55:@5176.4]
  wire [3:0] _T_5795; // @[Bitwise.scala 48:55:@5176.4]
  wire [1:0] _T_5796; // @[Bitwise.scala 48:55:@5177.4]
  wire [1:0] _GEN_807; // @[Bitwise.scala 48:55:@5178.4]
  wire [2:0] _T_5797; // @[Bitwise.scala 48:55:@5178.4]
  wire [1:0] _T_5798; // @[Bitwise.scala 48:55:@5179.4]
  wire [1:0] _GEN_808; // @[Bitwise.scala 48:55:@5180.4]
  wire [2:0] _T_5799; // @[Bitwise.scala 48:55:@5180.4]
  wire [3:0] _T_5800; // @[Bitwise.scala 48:55:@5181.4]
  wire [4:0] _T_5801; // @[Bitwise.scala 48:55:@5182.4]
  wire [1:0] _T_5802; // @[Bitwise.scala 48:55:@5183.4]
  wire [1:0] _T_5803; // @[Bitwise.scala 48:55:@5184.4]
  wire [1:0] _GEN_809; // @[Bitwise.scala 48:55:@5185.4]
  wire [2:0] _T_5804; // @[Bitwise.scala 48:55:@5185.4]
  wire [2:0] _GEN_810; // @[Bitwise.scala 48:55:@5186.4]
  wire [3:0] _T_5805; // @[Bitwise.scala 48:55:@5186.4]
  wire [1:0] _T_5806; // @[Bitwise.scala 48:55:@5187.4]
  wire [1:0] _GEN_811; // @[Bitwise.scala 48:55:@5188.4]
  wire [2:0] _T_5807; // @[Bitwise.scala 48:55:@5188.4]
  wire [1:0] _T_5808; // @[Bitwise.scala 48:55:@5189.4]
  wire [1:0] _GEN_812; // @[Bitwise.scala 48:55:@5190.4]
  wire [2:0] _T_5809; // @[Bitwise.scala 48:55:@5190.4]
  wire [3:0] _T_5810; // @[Bitwise.scala 48:55:@5191.4]
  wire [4:0] _T_5811; // @[Bitwise.scala 48:55:@5192.4]
  wire [5:0] _T_5812; // @[Bitwise.scala 48:55:@5193.4]
  wire [6:0] _T_5813; // @[Bitwise.scala 48:55:@5194.4]
  wire [44:0] _T_5877; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5259.4]
  wire  _T_5878; // @[Bitwise.scala 50:65:@5260.4]
  wire  _T_5879; // @[Bitwise.scala 50:65:@5261.4]
  wire  _T_5880; // @[Bitwise.scala 50:65:@5262.4]
  wire  _T_5881; // @[Bitwise.scala 50:65:@5263.4]
  wire  _T_5882; // @[Bitwise.scala 50:65:@5264.4]
  wire  _T_5883; // @[Bitwise.scala 50:65:@5265.4]
  wire  _T_5884; // @[Bitwise.scala 50:65:@5266.4]
  wire  _T_5885; // @[Bitwise.scala 50:65:@5267.4]
  wire  _T_5886; // @[Bitwise.scala 50:65:@5268.4]
  wire  _T_5887; // @[Bitwise.scala 50:65:@5269.4]
  wire  _T_5888; // @[Bitwise.scala 50:65:@5270.4]
  wire  _T_5889; // @[Bitwise.scala 50:65:@5271.4]
  wire  _T_5890; // @[Bitwise.scala 50:65:@5272.4]
  wire  _T_5891; // @[Bitwise.scala 50:65:@5273.4]
  wire  _T_5892; // @[Bitwise.scala 50:65:@5274.4]
  wire  _T_5893; // @[Bitwise.scala 50:65:@5275.4]
  wire  _T_5894; // @[Bitwise.scala 50:65:@5276.4]
  wire  _T_5895; // @[Bitwise.scala 50:65:@5277.4]
  wire  _T_5896; // @[Bitwise.scala 50:65:@5278.4]
  wire  _T_5897; // @[Bitwise.scala 50:65:@5279.4]
  wire  _T_5898; // @[Bitwise.scala 50:65:@5280.4]
  wire  _T_5899; // @[Bitwise.scala 50:65:@5281.4]
  wire  _T_5900; // @[Bitwise.scala 50:65:@5282.4]
  wire  _T_5901; // @[Bitwise.scala 50:65:@5283.4]
  wire  _T_5902; // @[Bitwise.scala 50:65:@5284.4]
  wire  _T_5903; // @[Bitwise.scala 50:65:@5285.4]
  wire  _T_5904; // @[Bitwise.scala 50:65:@5286.4]
  wire  _T_5905; // @[Bitwise.scala 50:65:@5287.4]
  wire  _T_5906; // @[Bitwise.scala 50:65:@5288.4]
  wire  _T_5907; // @[Bitwise.scala 50:65:@5289.4]
  wire  _T_5908; // @[Bitwise.scala 50:65:@5290.4]
  wire  _T_5909; // @[Bitwise.scala 50:65:@5291.4]
  wire  _T_5910; // @[Bitwise.scala 50:65:@5292.4]
  wire  _T_5911; // @[Bitwise.scala 50:65:@5293.4]
  wire  _T_5912; // @[Bitwise.scala 50:65:@5294.4]
  wire  _T_5913; // @[Bitwise.scala 50:65:@5295.4]
  wire  _T_5914; // @[Bitwise.scala 50:65:@5296.4]
  wire  _T_5915; // @[Bitwise.scala 50:65:@5297.4]
  wire  _T_5916; // @[Bitwise.scala 50:65:@5298.4]
  wire  _T_5917; // @[Bitwise.scala 50:65:@5299.4]
  wire  _T_5918; // @[Bitwise.scala 50:65:@5300.4]
  wire  _T_5919; // @[Bitwise.scala 50:65:@5301.4]
  wire  _T_5920; // @[Bitwise.scala 50:65:@5302.4]
  wire  _T_5921; // @[Bitwise.scala 50:65:@5303.4]
  wire  _T_5922; // @[Bitwise.scala 50:65:@5304.4]
  wire [1:0] _T_5923; // @[Bitwise.scala 48:55:@5305.4]
  wire [1:0] _T_5924; // @[Bitwise.scala 48:55:@5306.4]
  wire [1:0] _GEN_813; // @[Bitwise.scala 48:55:@5307.4]
  wire [2:0] _T_5925; // @[Bitwise.scala 48:55:@5307.4]
  wire [2:0] _GEN_814; // @[Bitwise.scala 48:55:@5308.4]
  wire [3:0] _T_5926; // @[Bitwise.scala 48:55:@5308.4]
  wire [1:0] _T_5927; // @[Bitwise.scala 48:55:@5309.4]
  wire [1:0] _GEN_815; // @[Bitwise.scala 48:55:@5310.4]
  wire [2:0] _T_5928; // @[Bitwise.scala 48:55:@5310.4]
  wire [1:0] _T_5929; // @[Bitwise.scala 48:55:@5311.4]
  wire [1:0] _GEN_816; // @[Bitwise.scala 48:55:@5312.4]
  wire [2:0] _T_5930; // @[Bitwise.scala 48:55:@5312.4]
  wire [3:0] _T_5931; // @[Bitwise.scala 48:55:@5313.4]
  wire [4:0] _T_5932; // @[Bitwise.scala 48:55:@5314.4]
  wire [1:0] _T_5933; // @[Bitwise.scala 48:55:@5315.4]
  wire [1:0] _T_5934; // @[Bitwise.scala 48:55:@5316.4]
  wire [1:0] _GEN_817; // @[Bitwise.scala 48:55:@5317.4]
  wire [2:0] _T_5935; // @[Bitwise.scala 48:55:@5317.4]
  wire [2:0] _GEN_818; // @[Bitwise.scala 48:55:@5318.4]
  wire [3:0] _T_5936; // @[Bitwise.scala 48:55:@5318.4]
  wire [1:0] _T_5937; // @[Bitwise.scala 48:55:@5319.4]
  wire [1:0] _GEN_819; // @[Bitwise.scala 48:55:@5320.4]
  wire [2:0] _T_5938; // @[Bitwise.scala 48:55:@5320.4]
  wire [1:0] _T_5939; // @[Bitwise.scala 48:55:@5321.4]
  wire [1:0] _GEN_820; // @[Bitwise.scala 48:55:@5322.4]
  wire [2:0] _T_5940; // @[Bitwise.scala 48:55:@5322.4]
  wire [3:0] _T_5941; // @[Bitwise.scala 48:55:@5323.4]
  wire [4:0] _T_5942; // @[Bitwise.scala 48:55:@5324.4]
  wire [5:0] _T_5943; // @[Bitwise.scala 48:55:@5325.4]
  wire [1:0] _T_5944; // @[Bitwise.scala 48:55:@5326.4]
  wire [1:0] _T_5945; // @[Bitwise.scala 48:55:@5327.4]
  wire [1:0] _GEN_821; // @[Bitwise.scala 48:55:@5328.4]
  wire [2:0] _T_5946; // @[Bitwise.scala 48:55:@5328.4]
  wire [2:0] _GEN_822; // @[Bitwise.scala 48:55:@5329.4]
  wire [3:0] _T_5947; // @[Bitwise.scala 48:55:@5329.4]
  wire [1:0] _T_5948; // @[Bitwise.scala 48:55:@5330.4]
  wire [1:0] _GEN_823; // @[Bitwise.scala 48:55:@5331.4]
  wire [2:0] _T_5949; // @[Bitwise.scala 48:55:@5331.4]
  wire [1:0] _T_5950; // @[Bitwise.scala 48:55:@5332.4]
  wire [1:0] _GEN_824; // @[Bitwise.scala 48:55:@5333.4]
  wire [2:0] _T_5951; // @[Bitwise.scala 48:55:@5333.4]
  wire [3:0] _T_5952; // @[Bitwise.scala 48:55:@5334.4]
  wire [4:0] _T_5953; // @[Bitwise.scala 48:55:@5335.4]
  wire [1:0] _T_5954; // @[Bitwise.scala 48:55:@5336.4]
  wire [1:0] _GEN_825; // @[Bitwise.scala 48:55:@5337.4]
  wire [2:0] _T_5955; // @[Bitwise.scala 48:55:@5337.4]
  wire [1:0] _T_5956; // @[Bitwise.scala 48:55:@5338.4]
  wire [1:0] _GEN_826; // @[Bitwise.scala 48:55:@5339.4]
  wire [2:0] _T_5957; // @[Bitwise.scala 48:55:@5339.4]
  wire [3:0] _T_5958; // @[Bitwise.scala 48:55:@5340.4]
  wire [1:0] _T_5959; // @[Bitwise.scala 48:55:@5341.4]
  wire [1:0] _GEN_827; // @[Bitwise.scala 48:55:@5342.4]
  wire [2:0] _T_5960; // @[Bitwise.scala 48:55:@5342.4]
  wire [1:0] _T_5961; // @[Bitwise.scala 48:55:@5343.4]
  wire [1:0] _GEN_828; // @[Bitwise.scala 48:55:@5344.4]
  wire [2:0] _T_5962; // @[Bitwise.scala 48:55:@5344.4]
  wire [3:0] _T_5963; // @[Bitwise.scala 48:55:@5345.4]
  wire [4:0] _T_5964; // @[Bitwise.scala 48:55:@5346.4]
  wire [5:0] _T_5965; // @[Bitwise.scala 48:55:@5347.4]
  wire [6:0] _T_5966; // @[Bitwise.scala 48:55:@5348.4]
  wire [45:0] _T_6030; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5413.4]
  wire  _T_6031; // @[Bitwise.scala 50:65:@5414.4]
  wire  _T_6032; // @[Bitwise.scala 50:65:@5415.4]
  wire  _T_6033; // @[Bitwise.scala 50:65:@5416.4]
  wire  _T_6034; // @[Bitwise.scala 50:65:@5417.4]
  wire  _T_6035; // @[Bitwise.scala 50:65:@5418.4]
  wire  _T_6036; // @[Bitwise.scala 50:65:@5419.4]
  wire  _T_6037; // @[Bitwise.scala 50:65:@5420.4]
  wire  _T_6038; // @[Bitwise.scala 50:65:@5421.4]
  wire  _T_6039; // @[Bitwise.scala 50:65:@5422.4]
  wire  _T_6040; // @[Bitwise.scala 50:65:@5423.4]
  wire  _T_6041; // @[Bitwise.scala 50:65:@5424.4]
  wire  _T_6042; // @[Bitwise.scala 50:65:@5425.4]
  wire  _T_6043; // @[Bitwise.scala 50:65:@5426.4]
  wire  _T_6044; // @[Bitwise.scala 50:65:@5427.4]
  wire  _T_6045; // @[Bitwise.scala 50:65:@5428.4]
  wire  _T_6046; // @[Bitwise.scala 50:65:@5429.4]
  wire  _T_6047; // @[Bitwise.scala 50:65:@5430.4]
  wire  _T_6048; // @[Bitwise.scala 50:65:@5431.4]
  wire  _T_6049; // @[Bitwise.scala 50:65:@5432.4]
  wire  _T_6050; // @[Bitwise.scala 50:65:@5433.4]
  wire  _T_6051; // @[Bitwise.scala 50:65:@5434.4]
  wire  _T_6052; // @[Bitwise.scala 50:65:@5435.4]
  wire  _T_6053; // @[Bitwise.scala 50:65:@5436.4]
  wire  _T_6054; // @[Bitwise.scala 50:65:@5437.4]
  wire  _T_6055; // @[Bitwise.scala 50:65:@5438.4]
  wire  _T_6056; // @[Bitwise.scala 50:65:@5439.4]
  wire  _T_6057; // @[Bitwise.scala 50:65:@5440.4]
  wire  _T_6058; // @[Bitwise.scala 50:65:@5441.4]
  wire  _T_6059; // @[Bitwise.scala 50:65:@5442.4]
  wire  _T_6060; // @[Bitwise.scala 50:65:@5443.4]
  wire  _T_6061; // @[Bitwise.scala 50:65:@5444.4]
  wire  _T_6062; // @[Bitwise.scala 50:65:@5445.4]
  wire  _T_6063; // @[Bitwise.scala 50:65:@5446.4]
  wire  _T_6064; // @[Bitwise.scala 50:65:@5447.4]
  wire  _T_6065; // @[Bitwise.scala 50:65:@5448.4]
  wire  _T_6066; // @[Bitwise.scala 50:65:@5449.4]
  wire  _T_6067; // @[Bitwise.scala 50:65:@5450.4]
  wire  _T_6068; // @[Bitwise.scala 50:65:@5451.4]
  wire  _T_6069; // @[Bitwise.scala 50:65:@5452.4]
  wire  _T_6070; // @[Bitwise.scala 50:65:@5453.4]
  wire  _T_6071; // @[Bitwise.scala 50:65:@5454.4]
  wire  _T_6072; // @[Bitwise.scala 50:65:@5455.4]
  wire  _T_6073; // @[Bitwise.scala 50:65:@5456.4]
  wire  _T_6074; // @[Bitwise.scala 50:65:@5457.4]
  wire  _T_6075; // @[Bitwise.scala 50:65:@5458.4]
  wire  _T_6076; // @[Bitwise.scala 50:65:@5459.4]
  wire [1:0] _T_6077; // @[Bitwise.scala 48:55:@5460.4]
  wire [1:0] _T_6078; // @[Bitwise.scala 48:55:@5461.4]
  wire [1:0] _GEN_829; // @[Bitwise.scala 48:55:@5462.4]
  wire [2:0] _T_6079; // @[Bitwise.scala 48:55:@5462.4]
  wire [2:0] _GEN_830; // @[Bitwise.scala 48:55:@5463.4]
  wire [3:0] _T_6080; // @[Bitwise.scala 48:55:@5463.4]
  wire [1:0] _T_6081; // @[Bitwise.scala 48:55:@5464.4]
  wire [1:0] _GEN_831; // @[Bitwise.scala 48:55:@5465.4]
  wire [2:0] _T_6082; // @[Bitwise.scala 48:55:@5465.4]
  wire [1:0] _T_6083; // @[Bitwise.scala 48:55:@5466.4]
  wire [1:0] _GEN_832; // @[Bitwise.scala 48:55:@5467.4]
  wire [2:0] _T_6084; // @[Bitwise.scala 48:55:@5467.4]
  wire [3:0] _T_6085; // @[Bitwise.scala 48:55:@5468.4]
  wire [4:0] _T_6086; // @[Bitwise.scala 48:55:@5469.4]
  wire [1:0] _T_6087; // @[Bitwise.scala 48:55:@5470.4]
  wire [1:0] _GEN_833; // @[Bitwise.scala 48:55:@5471.4]
  wire [2:0] _T_6088; // @[Bitwise.scala 48:55:@5471.4]
  wire [1:0] _T_6089; // @[Bitwise.scala 48:55:@5472.4]
  wire [1:0] _GEN_834; // @[Bitwise.scala 48:55:@5473.4]
  wire [2:0] _T_6090; // @[Bitwise.scala 48:55:@5473.4]
  wire [3:0] _T_6091; // @[Bitwise.scala 48:55:@5474.4]
  wire [1:0] _T_6092; // @[Bitwise.scala 48:55:@5475.4]
  wire [1:0] _GEN_835; // @[Bitwise.scala 48:55:@5476.4]
  wire [2:0] _T_6093; // @[Bitwise.scala 48:55:@5476.4]
  wire [1:0] _T_6094; // @[Bitwise.scala 48:55:@5477.4]
  wire [1:0] _GEN_836; // @[Bitwise.scala 48:55:@5478.4]
  wire [2:0] _T_6095; // @[Bitwise.scala 48:55:@5478.4]
  wire [3:0] _T_6096; // @[Bitwise.scala 48:55:@5479.4]
  wire [4:0] _T_6097; // @[Bitwise.scala 48:55:@5480.4]
  wire [5:0] _T_6098; // @[Bitwise.scala 48:55:@5481.4]
  wire [1:0] _T_6099; // @[Bitwise.scala 48:55:@5482.4]
  wire [1:0] _T_6100; // @[Bitwise.scala 48:55:@5483.4]
  wire [1:0] _GEN_837; // @[Bitwise.scala 48:55:@5484.4]
  wire [2:0] _T_6101; // @[Bitwise.scala 48:55:@5484.4]
  wire [2:0] _GEN_838; // @[Bitwise.scala 48:55:@5485.4]
  wire [3:0] _T_6102; // @[Bitwise.scala 48:55:@5485.4]
  wire [1:0] _T_6103; // @[Bitwise.scala 48:55:@5486.4]
  wire [1:0] _GEN_839; // @[Bitwise.scala 48:55:@5487.4]
  wire [2:0] _T_6104; // @[Bitwise.scala 48:55:@5487.4]
  wire [1:0] _T_6105; // @[Bitwise.scala 48:55:@5488.4]
  wire [1:0] _GEN_840; // @[Bitwise.scala 48:55:@5489.4]
  wire [2:0] _T_6106; // @[Bitwise.scala 48:55:@5489.4]
  wire [3:0] _T_6107; // @[Bitwise.scala 48:55:@5490.4]
  wire [4:0] _T_6108; // @[Bitwise.scala 48:55:@5491.4]
  wire [1:0] _T_6109; // @[Bitwise.scala 48:55:@5492.4]
  wire [1:0] _GEN_841; // @[Bitwise.scala 48:55:@5493.4]
  wire [2:0] _T_6110; // @[Bitwise.scala 48:55:@5493.4]
  wire [1:0] _T_6111; // @[Bitwise.scala 48:55:@5494.4]
  wire [1:0] _GEN_842; // @[Bitwise.scala 48:55:@5495.4]
  wire [2:0] _T_6112; // @[Bitwise.scala 48:55:@5495.4]
  wire [3:0] _T_6113; // @[Bitwise.scala 48:55:@5496.4]
  wire [1:0] _T_6114; // @[Bitwise.scala 48:55:@5497.4]
  wire [1:0] _GEN_843; // @[Bitwise.scala 48:55:@5498.4]
  wire [2:0] _T_6115; // @[Bitwise.scala 48:55:@5498.4]
  wire [1:0] _T_6116; // @[Bitwise.scala 48:55:@5499.4]
  wire [1:0] _GEN_844; // @[Bitwise.scala 48:55:@5500.4]
  wire [2:0] _T_6117; // @[Bitwise.scala 48:55:@5500.4]
  wire [3:0] _T_6118; // @[Bitwise.scala 48:55:@5501.4]
  wire [4:0] _T_6119; // @[Bitwise.scala 48:55:@5502.4]
  wire [5:0] _T_6120; // @[Bitwise.scala 48:55:@5503.4]
  wire [6:0] _T_6121; // @[Bitwise.scala 48:55:@5504.4]
  wire [46:0] _T_6185; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5569.4]
  wire  _T_6186; // @[Bitwise.scala 50:65:@5570.4]
  wire  _T_6187; // @[Bitwise.scala 50:65:@5571.4]
  wire  _T_6188; // @[Bitwise.scala 50:65:@5572.4]
  wire  _T_6189; // @[Bitwise.scala 50:65:@5573.4]
  wire  _T_6190; // @[Bitwise.scala 50:65:@5574.4]
  wire  _T_6191; // @[Bitwise.scala 50:65:@5575.4]
  wire  _T_6192; // @[Bitwise.scala 50:65:@5576.4]
  wire  _T_6193; // @[Bitwise.scala 50:65:@5577.4]
  wire  _T_6194; // @[Bitwise.scala 50:65:@5578.4]
  wire  _T_6195; // @[Bitwise.scala 50:65:@5579.4]
  wire  _T_6196; // @[Bitwise.scala 50:65:@5580.4]
  wire  _T_6197; // @[Bitwise.scala 50:65:@5581.4]
  wire  _T_6198; // @[Bitwise.scala 50:65:@5582.4]
  wire  _T_6199; // @[Bitwise.scala 50:65:@5583.4]
  wire  _T_6200; // @[Bitwise.scala 50:65:@5584.4]
  wire  _T_6201; // @[Bitwise.scala 50:65:@5585.4]
  wire  _T_6202; // @[Bitwise.scala 50:65:@5586.4]
  wire  _T_6203; // @[Bitwise.scala 50:65:@5587.4]
  wire  _T_6204; // @[Bitwise.scala 50:65:@5588.4]
  wire  _T_6205; // @[Bitwise.scala 50:65:@5589.4]
  wire  _T_6206; // @[Bitwise.scala 50:65:@5590.4]
  wire  _T_6207; // @[Bitwise.scala 50:65:@5591.4]
  wire  _T_6208; // @[Bitwise.scala 50:65:@5592.4]
  wire  _T_6209; // @[Bitwise.scala 50:65:@5593.4]
  wire  _T_6210; // @[Bitwise.scala 50:65:@5594.4]
  wire  _T_6211; // @[Bitwise.scala 50:65:@5595.4]
  wire  _T_6212; // @[Bitwise.scala 50:65:@5596.4]
  wire  _T_6213; // @[Bitwise.scala 50:65:@5597.4]
  wire  _T_6214; // @[Bitwise.scala 50:65:@5598.4]
  wire  _T_6215; // @[Bitwise.scala 50:65:@5599.4]
  wire  _T_6216; // @[Bitwise.scala 50:65:@5600.4]
  wire  _T_6217; // @[Bitwise.scala 50:65:@5601.4]
  wire  _T_6218; // @[Bitwise.scala 50:65:@5602.4]
  wire  _T_6219; // @[Bitwise.scala 50:65:@5603.4]
  wire  _T_6220; // @[Bitwise.scala 50:65:@5604.4]
  wire  _T_6221; // @[Bitwise.scala 50:65:@5605.4]
  wire  _T_6222; // @[Bitwise.scala 50:65:@5606.4]
  wire  _T_6223; // @[Bitwise.scala 50:65:@5607.4]
  wire  _T_6224; // @[Bitwise.scala 50:65:@5608.4]
  wire  _T_6225; // @[Bitwise.scala 50:65:@5609.4]
  wire  _T_6226; // @[Bitwise.scala 50:65:@5610.4]
  wire  _T_6227; // @[Bitwise.scala 50:65:@5611.4]
  wire  _T_6228; // @[Bitwise.scala 50:65:@5612.4]
  wire  _T_6229; // @[Bitwise.scala 50:65:@5613.4]
  wire  _T_6230; // @[Bitwise.scala 50:65:@5614.4]
  wire  _T_6231; // @[Bitwise.scala 50:65:@5615.4]
  wire  _T_6232; // @[Bitwise.scala 50:65:@5616.4]
  wire [1:0] _T_6233; // @[Bitwise.scala 48:55:@5617.4]
  wire [1:0] _T_6234; // @[Bitwise.scala 48:55:@5618.4]
  wire [1:0] _GEN_845; // @[Bitwise.scala 48:55:@5619.4]
  wire [2:0] _T_6235; // @[Bitwise.scala 48:55:@5619.4]
  wire [2:0] _GEN_846; // @[Bitwise.scala 48:55:@5620.4]
  wire [3:0] _T_6236; // @[Bitwise.scala 48:55:@5620.4]
  wire [1:0] _T_6237; // @[Bitwise.scala 48:55:@5621.4]
  wire [1:0] _GEN_847; // @[Bitwise.scala 48:55:@5622.4]
  wire [2:0] _T_6238; // @[Bitwise.scala 48:55:@5622.4]
  wire [1:0] _T_6239; // @[Bitwise.scala 48:55:@5623.4]
  wire [1:0] _GEN_848; // @[Bitwise.scala 48:55:@5624.4]
  wire [2:0] _T_6240; // @[Bitwise.scala 48:55:@5624.4]
  wire [3:0] _T_6241; // @[Bitwise.scala 48:55:@5625.4]
  wire [4:0] _T_6242; // @[Bitwise.scala 48:55:@5626.4]
  wire [1:0] _T_6243; // @[Bitwise.scala 48:55:@5627.4]
  wire [1:0] _GEN_849; // @[Bitwise.scala 48:55:@5628.4]
  wire [2:0] _T_6244; // @[Bitwise.scala 48:55:@5628.4]
  wire [1:0] _T_6245; // @[Bitwise.scala 48:55:@5629.4]
  wire [1:0] _GEN_850; // @[Bitwise.scala 48:55:@5630.4]
  wire [2:0] _T_6246; // @[Bitwise.scala 48:55:@5630.4]
  wire [3:0] _T_6247; // @[Bitwise.scala 48:55:@5631.4]
  wire [1:0] _T_6248; // @[Bitwise.scala 48:55:@5632.4]
  wire [1:0] _GEN_851; // @[Bitwise.scala 48:55:@5633.4]
  wire [2:0] _T_6249; // @[Bitwise.scala 48:55:@5633.4]
  wire [1:0] _T_6250; // @[Bitwise.scala 48:55:@5634.4]
  wire [1:0] _GEN_852; // @[Bitwise.scala 48:55:@5635.4]
  wire [2:0] _T_6251; // @[Bitwise.scala 48:55:@5635.4]
  wire [3:0] _T_6252; // @[Bitwise.scala 48:55:@5636.4]
  wire [4:0] _T_6253; // @[Bitwise.scala 48:55:@5637.4]
  wire [5:0] _T_6254; // @[Bitwise.scala 48:55:@5638.4]
  wire [1:0] _T_6255; // @[Bitwise.scala 48:55:@5639.4]
  wire [1:0] _GEN_853; // @[Bitwise.scala 48:55:@5640.4]
  wire [2:0] _T_6256; // @[Bitwise.scala 48:55:@5640.4]
  wire [1:0] _T_6257; // @[Bitwise.scala 48:55:@5641.4]
  wire [1:0] _GEN_854; // @[Bitwise.scala 48:55:@5642.4]
  wire [2:0] _T_6258; // @[Bitwise.scala 48:55:@5642.4]
  wire [3:0] _T_6259; // @[Bitwise.scala 48:55:@5643.4]
  wire [1:0] _T_6260; // @[Bitwise.scala 48:55:@5644.4]
  wire [1:0] _GEN_855; // @[Bitwise.scala 48:55:@5645.4]
  wire [2:0] _T_6261; // @[Bitwise.scala 48:55:@5645.4]
  wire [1:0] _T_6262; // @[Bitwise.scala 48:55:@5646.4]
  wire [1:0] _GEN_856; // @[Bitwise.scala 48:55:@5647.4]
  wire [2:0] _T_6263; // @[Bitwise.scala 48:55:@5647.4]
  wire [3:0] _T_6264; // @[Bitwise.scala 48:55:@5648.4]
  wire [4:0] _T_6265; // @[Bitwise.scala 48:55:@5649.4]
  wire [1:0] _T_6266; // @[Bitwise.scala 48:55:@5650.4]
  wire [1:0] _GEN_857; // @[Bitwise.scala 48:55:@5651.4]
  wire [2:0] _T_6267; // @[Bitwise.scala 48:55:@5651.4]
  wire [1:0] _T_6268; // @[Bitwise.scala 48:55:@5652.4]
  wire [1:0] _GEN_858; // @[Bitwise.scala 48:55:@5653.4]
  wire [2:0] _T_6269; // @[Bitwise.scala 48:55:@5653.4]
  wire [3:0] _T_6270; // @[Bitwise.scala 48:55:@5654.4]
  wire [1:0] _T_6271; // @[Bitwise.scala 48:55:@5655.4]
  wire [1:0] _GEN_859; // @[Bitwise.scala 48:55:@5656.4]
  wire [2:0] _T_6272; // @[Bitwise.scala 48:55:@5656.4]
  wire [1:0] _T_6273; // @[Bitwise.scala 48:55:@5657.4]
  wire [1:0] _GEN_860; // @[Bitwise.scala 48:55:@5658.4]
  wire [2:0] _T_6274; // @[Bitwise.scala 48:55:@5658.4]
  wire [3:0] _T_6275; // @[Bitwise.scala 48:55:@5659.4]
  wire [4:0] _T_6276; // @[Bitwise.scala 48:55:@5660.4]
  wire [5:0] _T_6277; // @[Bitwise.scala 48:55:@5661.4]
  wire [6:0] _T_6278; // @[Bitwise.scala 48:55:@5662.4]
  wire [47:0] _T_6342; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5727.4]
  wire  _T_6343; // @[Bitwise.scala 50:65:@5728.4]
  wire  _T_6344; // @[Bitwise.scala 50:65:@5729.4]
  wire  _T_6345; // @[Bitwise.scala 50:65:@5730.4]
  wire  _T_6346; // @[Bitwise.scala 50:65:@5731.4]
  wire  _T_6347; // @[Bitwise.scala 50:65:@5732.4]
  wire  _T_6348; // @[Bitwise.scala 50:65:@5733.4]
  wire  _T_6349; // @[Bitwise.scala 50:65:@5734.4]
  wire  _T_6350; // @[Bitwise.scala 50:65:@5735.4]
  wire  _T_6351; // @[Bitwise.scala 50:65:@5736.4]
  wire  _T_6352; // @[Bitwise.scala 50:65:@5737.4]
  wire  _T_6353; // @[Bitwise.scala 50:65:@5738.4]
  wire  _T_6354; // @[Bitwise.scala 50:65:@5739.4]
  wire  _T_6355; // @[Bitwise.scala 50:65:@5740.4]
  wire  _T_6356; // @[Bitwise.scala 50:65:@5741.4]
  wire  _T_6357; // @[Bitwise.scala 50:65:@5742.4]
  wire  _T_6358; // @[Bitwise.scala 50:65:@5743.4]
  wire  _T_6359; // @[Bitwise.scala 50:65:@5744.4]
  wire  _T_6360; // @[Bitwise.scala 50:65:@5745.4]
  wire  _T_6361; // @[Bitwise.scala 50:65:@5746.4]
  wire  _T_6362; // @[Bitwise.scala 50:65:@5747.4]
  wire  _T_6363; // @[Bitwise.scala 50:65:@5748.4]
  wire  _T_6364; // @[Bitwise.scala 50:65:@5749.4]
  wire  _T_6365; // @[Bitwise.scala 50:65:@5750.4]
  wire  _T_6366; // @[Bitwise.scala 50:65:@5751.4]
  wire  _T_6367; // @[Bitwise.scala 50:65:@5752.4]
  wire  _T_6368; // @[Bitwise.scala 50:65:@5753.4]
  wire  _T_6369; // @[Bitwise.scala 50:65:@5754.4]
  wire  _T_6370; // @[Bitwise.scala 50:65:@5755.4]
  wire  _T_6371; // @[Bitwise.scala 50:65:@5756.4]
  wire  _T_6372; // @[Bitwise.scala 50:65:@5757.4]
  wire  _T_6373; // @[Bitwise.scala 50:65:@5758.4]
  wire  _T_6374; // @[Bitwise.scala 50:65:@5759.4]
  wire  _T_6375; // @[Bitwise.scala 50:65:@5760.4]
  wire  _T_6376; // @[Bitwise.scala 50:65:@5761.4]
  wire  _T_6377; // @[Bitwise.scala 50:65:@5762.4]
  wire  _T_6378; // @[Bitwise.scala 50:65:@5763.4]
  wire  _T_6379; // @[Bitwise.scala 50:65:@5764.4]
  wire  _T_6380; // @[Bitwise.scala 50:65:@5765.4]
  wire  _T_6381; // @[Bitwise.scala 50:65:@5766.4]
  wire  _T_6382; // @[Bitwise.scala 50:65:@5767.4]
  wire  _T_6383; // @[Bitwise.scala 50:65:@5768.4]
  wire  _T_6384; // @[Bitwise.scala 50:65:@5769.4]
  wire  _T_6385; // @[Bitwise.scala 50:65:@5770.4]
  wire  _T_6386; // @[Bitwise.scala 50:65:@5771.4]
  wire  _T_6387; // @[Bitwise.scala 50:65:@5772.4]
  wire  _T_6388; // @[Bitwise.scala 50:65:@5773.4]
  wire  _T_6389; // @[Bitwise.scala 50:65:@5774.4]
  wire  _T_6390; // @[Bitwise.scala 50:65:@5775.4]
  wire [1:0] _T_6391; // @[Bitwise.scala 48:55:@5776.4]
  wire [1:0] _GEN_861; // @[Bitwise.scala 48:55:@5777.4]
  wire [2:0] _T_6392; // @[Bitwise.scala 48:55:@5777.4]
  wire [1:0] _T_6393; // @[Bitwise.scala 48:55:@5778.4]
  wire [1:0] _GEN_862; // @[Bitwise.scala 48:55:@5779.4]
  wire [2:0] _T_6394; // @[Bitwise.scala 48:55:@5779.4]
  wire [3:0] _T_6395; // @[Bitwise.scala 48:55:@5780.4]
  wire [1:0] _T_6396; // @[Bitwise.scala 48:55:@5781.4]
  wire [1:0] _GEN_863; // @[Bitwise.scala 48:55:@5782.4]
  wire [2:0] _T_6397; // @[Bitwise.scala 48:55:@5782.4]
  wire [1:0] _T_6398; // @[Bitwise.scala 48:55:@5783.4]
  wire [1:0] _GEN_864; // @[Bitwise.scala 48:55:@5784.4]
  wire [2:0] _T_6399; // @[Bitwise.scala 48:55:@5784.4]
  wire [3:0] _T_6400; // @[Bitwise.scala 48:55:@5785.4]
  wire [4:0] _T_6401; // @[Bitwise.scala 48:55:@5786.4]
  wire [1:0] _T_6402; // @[Bitwise.scala 48:55:@5787.4]
  wire [1:0] _GEN_865; // @[Bitwise.scala 48:55:@5788.4]
  wire [2:0] _T_6403; // @[Bitwise.scala 48:55:@5788.4]
  wire [1:0] _T_6404; // @[Bitwise.scala 48:55:@5789.4]
  wire [1:0] _GEN_866; // @[Bitwise.scala 48:55:@5790.4]
  wire [2:0] _T_6405; // @[Bitwise.scala 48:55:@5790.4]
  wire [3:0] _T_6406; // @[Bitwise.scala 48:55:@5791.4]
  wire [1:0] _T_6407; // @[Bitwise.scala 48:55:@5792.4]
  wire [1:0] _GEN_867; // @[Bitwise.scala 48:55:@5793.4]
  wire [2:0] _T_6408; // @[Bitwise.scala 48:55:@5793.4]
  wire [1:0] _T_6409; // @[Bitwise.scala 48:55:@5794.4]
  wire [1:0] _GEN_868; // @[Bitwise.scala 48:55:@5795.4]
  wire [2:0] _T_6410; // @[Bitwise.scala 48:55:@5795.4]
  wire [3:0] _T_6411; // @[Bitwise.scala 48:55:@5796.4]
  wire [4:0] _T_6412; // @[Bitwise.scala 48:55:@5797.4]
  wire [5:0] _T_6413; // @[Bitwise.scala 48:55:@5798.4]
  wire [1:0] _T_6414; // @[Bitwise.scala 48:55:@5799.4]
  wire [1:0] _GEN_869; // @[Bitwise.scala 48:55:@5800.4]
  wire [2:0] _T_6415; // @[Bitwise.scala 48:55:@5800.4]
  wire [1:0] _T_6416; // @[Bitwise.scala 48:55:@5801.4]
  wire [1:0] _GEN_870; // @[Bitwise.scala 48:55:@5802.4]
  wire [2:0] _T_6417; // @[Bitwise.scala 48:55:@5802.4]
  wire [3:0] _T_6418; // @[Bitwise.scala 48:55:@5803.4]
  wire [1:0] _T_6419; // @[Bitwise.scala 48:55:@5804.4]
  wire [1:0] _GEN_871; // @[Bitwise.scala 48:55:@5805.4]
  wire [2:0] _T_6420; // @[Bitwise.scala 48:55:@5805.4]
  wire [1:0] _T_6421; // @[Bitwise.scala 48:55:@5806.4]
  wire [1:0] _GEN_872; // @[Bitwise.scala 48:55:@5807.4]
  wire [2:0] _T_6422; // @[Bitwise.scala 48:55:@5807.4]
  wire [3:0] _T_6423; // @[Bitwise.scala 48:55:@5808.4]
  wire [4:0] _T_6424; // @[Bitwise.scala 48:55:@5809.4]
  wire [1:0] _T_6425; // @[Bitwise.scala 48:55:@5810.4]
  wire [1:0] _GEN_873; // @[Bitwise.scala 48:55:@5811.4]
  wire [2:0] _T_6426; // @[Bitwise.scala 48:55:@5811.4]
  wire [1:0] _T_6427; // @[Bitwise.scala 48:55:@5812.4]
  wire [1:0] _GEN_874; // @[Bitwise.scala 48:55:@5813.4]
  wire [2:0] _T_6428; // @[Bitwise.scala 48:55:@5813.4]
  wire [3:0] _T_6429; // @[Bitwise.scala 48:55:@5814.4]
  wire [1:0] _T_6430; // @[Bitwise.scala 48:55:@5815.4]
  wire [1:0] _GEN_875; // @[Bitwise.scala 48:55:@5816.4]
  wire [2:0] _T_6431; // @[Bitwise.scala 48:55:@5816.4]
  wire [1:0] _T_6432; // @[Bitwise.scala 48:55:@5817.4]
  wire [1:0] _GEN_876; // @[Bitwise.scala 48:55:@5818.4]
  wire [2:0] _T_6433; // @[Bitwise.scala 48:55:@5818.4]
  wire [3:0] _T_6434; // @[Bitwise.scala 48:55:@5819.4]
  wire [4:0] _T_6435; // @[Bitwise.scala 48:55:@5820.4]
  wire [5:0] _T_6436; // @[Bitwise.scala 48:55:@5821.4]
  wire [6:0] _T_6437; // @[Bitwise.scala 48:55:@5822.4]
  wire [48:0] _T_6501; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5887.4]
  wire  _T_6502; // @[Bitwise.scala 50:65:@5888.4]
  wire  _T_6503; // @[Bitwise.scala 50:65:@5889.4]
  wire  _T_6504; // @[Bitwise.scala 50:65:@5890.4]
  wire  _T_6505; // @[Bitwise.scala 50:65:@5891.4]
  wire  _T_6506; // @[Bitwise.scala 50:65:@5892.4]
  wire  _T_6507; // @[Bitwise.scala 50:65:@5893.4]
  wire  _T_6508; // @[Bitwise.scala 50:65:@5894.4]
  wire  _T_6509; // @[Bitwise.scala 50:65:@5895.4]
  wire  _T_6510; // @[Bitwise.scala 50:65:@5896.4]
  wire  _T_6511; // @[Bitwise.scala 50:65:@5897.4]
  wire  _T_6512; // @[Bitwise.scala 50:65:@5898.4]
  wire  _T_6513; // @[Bitwise.scala 50:65:@5899.4]
  wire  _T_6514; // @[Bitwise.scala 50:65:@5900.4]
  wire  _T_6515; // @[Bitwise.scala 50:65:@5901.4]
  wire  _T_6516; // @[Bitwise.scala 50:65:@5902.4]
  wire  _T_6517; // @[Bitwise.scala 50:65:@5903.4]
  wire  _T_6518; // @[Bitwise.scala 50:65:@5904.4]
  wire  _T_6519; // @[Bitwise.scala 50:65:@5905.4]
  wire  _T_6520; // @[Bitwise.scala 50:65:@5906.4]
  wire  _T_6521; // @[Bitwise.scala 50:65:@5907.4]
  wire  _T_6522; // @[Bitwise.scala 50:65:@5908.4]
  wire  _T_6523; // @[Bitwise.scala 50:65:@5909.4]
  wire  _T_6524; // @[Bitwise.scala 50:65:@5910.4]
  wire  _T_6525; // @[Bitwise.scala 50:65:@5911.4]
  wire  _T_6526; // @[Bitwise.scala 50:65:@5912.4]
  wire  _T_6527; // @[Bitwise.scala 50:65:@5913.4]
  wire  _T_6528; // @[Bitwise.scala 50:65:@5914.4]
  wire  _T_6529; // @[Bitwise.scala 50:65:@5915.4]
  wire  _T_6530; // @[Bitwise.scala 50:65:@5916.4]
  wire  _T_6531; // @[Bitwise.scala 50:65:@5917.4]
  wire  _T_6532; // @[Bitwise.scala 50:65:@5918.4]
  wire  _T_6533; // @[Bitwise.scala 50:65:@5919.4]
  wire  _T_6534; // @[Bitwise.scala 50:65:@5920.4]
  wire  _T_6535; // @[Bitwise.scala 50:65:@5921.4]
  wire  _T_6536; // @[Bitwise.scala 50:65:@5922.4]
  wire  _T_6537; // @[Bitwise.scala 50:65:@5923.4]
  wire  _T_6538; // @[Bitwise.scala 50:65:@5924.4]
  wire  _T_6539; // @[Bitwise.scala 50:65:@5925.4]
  wire  _T_6540; // @[Bitwise.scala 50:65:@5926.4]
  wire  _T_6541; // @[Bitwise.scala 50:65:@5927.4]
  wire  _T_6542; // @[Bitwise.scala 50:65:@5928.4]
  wire  _T_6543; // @[Bitwise.scala 50:65:@5929.4]
  wire  _T_6544; // @[Bitwise.scala 50:65:@5930.4]
  wire  _T_6545; // @[Bitwise.scala 50:65:@5931.4]
  wire  _T_6546; // @[Bitwise.scala 50:65:@5932.4]
  wire  _T_6547; // @[Bitwise.scala 50:65:@5933.4]
  wire  _T_6548; // @[Bitwise.scala 50:65:@5934.4]
  wire  _T_6549; // @[Bitwise.scala 50:65:@5935.4]
  wire  _T_6550; // @[Bitwise.scala 50:65:@5936.4]
  wire [1:0] _T_6551; // @[Bitwise.scala 48:55:@5937.4]
  wire [1:0] _GEN_877; // @[Bitwise.scala 48:55:@5938.4]
  wire [2:0] _T_6552; // @[Bitwise.scala 48:55:@5938.4]
  wire [1:0] _T_6553; // @[Bitwise.scala 48:55:@5939.4]
  wire [1:0] _GEN_878; // @[Bitwise.scala 48:55:@5940.4]
  wire [2:0] _T_6554; // @[Bitwise.scala 48:55:@5940.4]
  wire [3:0] _T_6555; // @[Bitwise.scala 48:55:@5941.4]
  wire [1:0] _T_6556; // @[Bitwise.scala 48:55:@5942.4]
  wire [1:0] _GEN_879; // @[Bitwise.scala 48:55:@5943.4]
  wire [2:0] _T_6557; // @[Bitwise.scala 48:55:@5943.4]
  wire [1:0] _T_6558; // @[Bitwise.scala 48:55:@5944.4]
  wire [1:0] _GEN_880; // @[Bitwise.scala 48:55:@5945.4]
  wire [2:0] _T_6559; // @[Bitwise.scala 48:55:@5945.4]
  wire [3:0] _T_6560; // @[Bitwise.scala 48:55:@5946.4]
  wire [4:0] _T_6561; // @[Bitwise.scala 48:55:@5947.4]
  wire [1:0] _T_6562; // @[Bitwise.scala 48:55:@5948.4]
  wire [1:0] _GEN_881; // @[Bitwise.scala 48:55:@5949.4]
  wire [2:0] _T_6563; // @[Bitwise.scala 48:55:@5949.4]
  wire [1:0] _T_6564; // @[Bitwise.scala 48:55:@5950.4]
  wire [1:0] _GEN_882; // @[Bitwise.scala 48:55:@5951.4]
  wire [2:0] _T_6565; // @[Bitwise.scala 48:55:@5951.4]
  wire [3:0] _T_6566; // @[Bitwise.scala 48:55:@5952.4]
  wire [1:0] _T_6567; // @[Bitwise.scala 48:55:@5953.4]
  wire [1:0] _GEN_883; // @[Bitwise.scala 48:55:@5954.4]
  wire [2:0] _T_6568; // @[Bitwise.scala 48:55:@5954.4]
  wire [1:0] _T_6569; // @[Bitwise.scala 48:55:@5955.4]
  wire [1:0] _GEN_884; // @[Bitwise.scala 48:55:@5956.4]
  wire [2:0] _T_6570; // @[Bitwise.scala 48:55:@5956.4]
  wire [3:0] _T_6571; // @[Bitwise.scala 48:55:@5957.4]
  wire [4:0] _T_6572; // @[Bitwise.scala 48:55:@5958.4]
  wire [5:0] _T_6573; // @[Bitwise.scala 48:55:@5959.4]
  wire [1:0] _T_6574; // @[Bitwise.scala 48:55:@5960.4]
  wire [1:0] _GEN_885; // @[Bitwise.scala 48:55:@5961.4]
  wire [2:0] _T_6575; // @[Bitwise.scala 48:55:@5961.4]
  wire [1:0] _T_6576; // @[Bitwise.scala 48:55:@5962.4]
  wire [1:0] _GEN_886; // @[Bitwise.scala 48:55:@5963.4]
  wire [2:0] _T_6577; // @[Bitwise.scala 48:55:@5963.4]
  wire [3:0] _T_6578; // @[Bitwise.scala 48:55:@5964.4]
  wire [1:0] _T_6579; // @[Bitwise.scala 48:55:@5965.4]
  wire [1:0] _GEN_887; // @[Bitwise.scala 48:55:@5966.4]
  wire [2:0] _T_6580; // @[Bitwise.scala 48:55:@5966.4]
  wire [1:0] _T_6581; // @[Bitwise.scala 48:55:@5967.4]
  wire [1:0] _GEN_888; // @[Bitwise.scala 48:55:@5968.4]
  wire [2:0] _T_6582; // @[Bitwise.scala 48:55:@5968.4]
  wire [3:0] _T_6583; // @[Bitwise.scala 48:55:@5969.4]
  wire [4:0] _T_6584; // @[Bitwise.scala 48:55:@5970.4]
  wire [1:0] _T_6585; // @[Bitwise.scala 48:55:@5971.4]
  wire [1:0] _GEN_889; // @[Bitwise.scala 48:55:@5972.4]
  wire [2:0] _T_6586; // @[Bitwise.scala 48:55:@5972.4]
  wire [1:0] _T_6587; // @[Bitwise.scala 48:55:@5973.4]
  wire [1:0] _GEN_890; // @[Bitwise.scala 48:55:@5974.4]
  wire [2:0] _T_6588; // @[Bitwise.scala 48:55:@5974.4]
  wire [3:0] _T_6589; // @[Bitwise.scala 48:55:@5975.4]
  wire [1:0] _T_6590; // @[Bitwise.scala 48:55:@5976.4]
  wire [1:0] _GEN_891; // @[Bitwise.scala 48:55:@5977.4]
  wire [2:0] _T_6591; // @[Bitwise.scala 48:55:@5977.4]
  wire [1:0] _T_6592; // @[Bitwise.scala 48:55:@5978.4]
  wire [1:0] _T_6593; // @[Bitwise.scala 48:55:@5979.4]
  wire [2:0] _T_6594; // @[Bitwise.scala 48:55:@5980.4]
  wire [3:0] _T_6595; // @[Bitwise.scala 48:55:@5981.4]
  wire [4:0] _T_6596; // @[Bitwise.scala 48:55:@5982.4]
  wire [5:0] _T_6597; // @[Bitwise.scala 48:55:@5983.4]
  wire [6:0] _T_6598; // @[Bitwise.scala 48:55:@5984.4]
  wire [49:0] _T_6662; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6049.4]
  wire  _T_6663; // @[Bitwise.scala 50:65:@6050.4]
  wire  _T_6664; // @[Bitwise.scala 50:65:@6051.4]
  wire  _T_6665; // @[Bitwise.scala 50:65:@6052.4]
  wire  _T_6666; // @[Bitwise.scala 50:65:@6053.4]
  wire  _T_6667; // @[Bitwise.scala 50:65:@6054.4]
  wire  _T_6668; // @[Bitwise.scala 50:65:@6055.4]
  wire  _T_6669; // @[Bitwise.scala 50:65:@6056.4]
  wire  _T_6670; // @[Bitwise.scala 50:65:@6057.4]
  wire  _T_6671; // @[Bitwise.scala 50:65:@6058.4]
  wire  _T_6672; // @[Bitwise.scala 50:65:@6059.4]
  wire  _T_6673; // @[Bitwise.scala 50:65:@6060.4]
  wire  _T_6674; // @[Bitwise.scala 50:65:@6061.4]
  wire  _T_6675; // @[Bitwise.scala 50:65:@6062.4]
  wire  _T_6676; // @[Bitwise.scala 50:65:@6063.4]
  wire  _T_6677; // @[Bitwise.scala 50:65:@6064.4]
  wire  _T_6678; // @[Bitwise.scala 50:65:@6065.4]
  wire  _T_6679; // @[Bitwise.scala 50:65:@6066.4]
  wire  _T_6680; // @[Bitwise.scala 50:65:@6067.4]
  wire  _T_6681; // @[Bitwise.scala 50:65:@6068.4]
  wire  _T_6682; // @[Bitwise.scala 50:65:@6069.4]
  wire  _T_6683; // @[Bitwise.scala 50:65:@6070.4]
  wire  _T_6684; // @[Bitwise.scala 50:65:@6071.4]
  wire  _T_6685; // @[Bitwise.scala 50:65:@6072.4]
  wire  _T_6686; // @[Bitwise.scala 50:65:@6073.4]
  wire  _T_6687; // @[Bitwise.scala 50:65:@6074.4]
  wire  _T_6688; // @[Bitwise.scala 50:65:@6075.4]
  wire  _T_6689; // @[Bitwise.scala 50:65:@6076.4]
  wire  _T_6690; // @[Bitwise.scala 50:65:@6077.4]
  wire  _T_6691; // @[Bitwise.scala 50:65:@6078.4]
  wire  _T_6692; // @[Bitwise.scala 50:65:@6079.4]
  wire  _T_6693; // @[Bitwise.scala 50:65:@6080.4]
  wire  _T_6694; // @[Bitwise.scala 50:65:@6081.4]
  wire  _T_6695; // @[Bitwise.scala 50:65:@6082.4]
  wire  _T_6696; // @[Bitwise.scala 50:65:@6083.4]
  wire  _T_6697; // @[Bitwise.scala 50:65:@6084.4]
  wire  _T_6698; // @[Bitwise.scala 50:65:@6085.4]
  wire  _T_6699; // @[Bitwise.scala 50:65:@6086.4]
  wire  _T_6700; // @[Bitwise.scala 50:65:@6087.4]
  wire  _T_6701; // @[Bitwise.scala 50:65:@6088.4]
  wire  _T_6702; // @[Bitwise.scala 50:65:@6089.4]
  wire  _T_6703; // @[Bitwise.scala 50:65:@6090.4]
  wire  _T_6704; // @[Bitwise.scala 50:65:@6091.4]
  wire  _T_6705; // @[Bitwise.scala 50:65:@6092.4]
  wire  _T_6706; // @[Bitwise.scala 50:65:@6093.4]
  wire  _T_6707; // @[Bitwise.scala 50:65:@6094.4]
  wire  _T_6708; // @[Bitwise.scala 50:65:@6095.4]
  wire  _T_6709; // @[Bitwise.scala 50:65:@6096.4]
  wire  _T_6710; // @[Bitwise.scala 50:65:@6097.4]
  wire  _T_6711; // @[Bitwise.scala 50:65:@6098.4]
  wire  _T_6712; // @[Bitwise.scala 50:65:@6099.4]
  wire [1:0] _T_6713; // @[Bitwise.scala 48:55:@6100.4]
  wire [1:0] _GEN_892; // @[Bitwise.scala 48:55:@6101.4]
  wire [2:0] _T_6714; // @[Bitwise.scala 48:55:@6101.4]
  wire [1:0] _T_6715; // @[Bitwise.scala 48:55:@6102.4]
  wire [1:0] _GEN_893; // @[Bitwise.scala 48:55:@6103.4]
  wire [2:0] _T_6716; // @[Bitwise.scala 48:55:@6103.4]
  wire [3:0] _T_6717; // @[Bitwise.scala 48:55:@6104.4]
  wire [1:0] _T_6718; // @[Bitwise.scala 48:55:@6105.4]
  wire [1:0] _GEN_894; // @[Bitwise.scala 48:55:@6106.4]
  wire [2:0] _T_6719; // @[Bitwise.scala 48:55:@6106.4]
  wire [1:0] _T_6720; // @[Bitwise.scala 48:55:@6107.4]
  wire [1:0] _GEN_895; // @[Bitwise.scala 48:55:@6108.4]
  wire [2:0] _T_6721; // @[Bitwise.scala 48:55:@6108.4]
  wire [3:0] _T_6722; // @[Bitwise.scala 48:55:@6109.4]
  wire [4:0] _T_6723; // @[Bitwise.scala 48:55:@6110.4]
  wire [1:0] _T_6724; // @[Bitwise.scala 48:55:@6111.4]
  wire [1:0] _GEN_896; // @[Bitwise.scala 48:55:@6112.4]
  wire [2:0] _T_6725; // @[Bitwise.scala 48:55:@6112.4]
  wire [1:0] _T_6726; // @[Bitwise.scala 48:55:@6113.4]
  wire [1:0] _GEN_897; // @[Bitwise.scala 48:55:@6114.4]
  wire [2:0] _T_6727; // @[Bitwise.scala 48:55:@6114.4]
  wire [3:0] _T_6728; // @[Bitwise.scala 48:55:@6115.4]
  wire [1:0] _T_6729; // @[Bitwise.scala 48:55:@6116.4]
  wire [1:0] _GEN_898; // @[Bitwise.scala 48:55:@6117.4]
  wire [2:0] _T_6730; // @[Bitwise.scala 48:55:@6117.4]
  wire [1:0] _T_6731; // @[Bitwise.scala 48:55:@6118.4]
  wire [1:0] _T_6732; // @[Bitwise.scala 48:55:@6119.4]
  wire [2:0] _T_6733; // @[Bitwise.scala 48:55:@6120.4]
  wire [3:0] _T_6734; // @[Bitwise.scala 48:55:@6121.4]
  wire [4:0] _T_6735; // @[Bitwise.scala 48:55:@6122.4]
  wire [5:0] _T_6736; // @[Bitwise.scala 48:55:@6123.4]
  wire [1:0] _T_6737; // @[Bitwise.scala 48:55:@6124.4]
  wire [1:0] _GEN_899; // @[Bitwise.scala 48:55:@6125.4]
  wire [2:0] _T_6738; // @[Bitwise.scala 48:55:@6125.4]
  wire [1:0] _T_6739; // @[Bitwise.scala 48:55:@6126.4]
  wire [1:0] _GEN_900; // @[Bitwise.scala 48:55:@6127.4]
  wire [2:0] _T_6740; // @[Bitwise.scala 48:55:@6127.4]
  wire [3:0] _T_6741; // @[Bitwise.scala 48:55:@6128.4]
  wire [1:0] _T_6742; // @[Bitwise.scala 48:55:@6129.4]
  wire [1:0] _GEN_901; // @[Bitwise.scala 48:55:@6130.4]
  wire [2:0] _T_6743; // @[Bitwise.scala 48:55:@6130.4]
  wire [1:0] _T_6744; // @[Bitwise.scala 48:55:@6131.4]
  wire [1:0] _GEN_902; // @[Bitwise.scala 48:55:@6132.4]
  wire [2:0] _T_6745; // @[Bitwise.scala 48:55:@6132.4]
  wire [3:0] _T_6746; // @[Bitwise.scala 48:55:@6133.4]
  wire [4:0] _T_6747; // @[Bitwise.scala 48:55:@6134.4]
  wire [1:0] _T_6748; // @[Bitwise.scala 48:55:@6135.4]
  wire [1:0] _GEN_903; // @[Bitwise.scala 48:55:@6136.4]
  wire [2:0] _T_6749; // @[Bitwise.scala 48:55:@6136.4]
  wire [1:0] _T_6750; // @[Bitwise.scala 48:55:@6137.4]
  wire [1:0] _GEN_904; // @[Bitwise.scala 48:55:@6138.4]
  wire [2:0] _T_6751; // @[Bitwise.scala 48:55:@6138.4]
  wire [3:0] _T_6752; // @[Bitwise.scala 48:55:@6139.4]
  wire [1:0] _T_6753; // @[Bitwise.scala 48:55:@6140.4]
  wire [1:0] _GEN_905; // @[Bitwise.scala 48:55:@6141.4]
  wire [2:0] _T_6754; // @[Bitwise.scala 48:55:@6141.4]
  wire [1:0] _T_6755; // @[Bitwise.scala 48:55:@6142.4]
  wire [1:0] _T_6756; // @[Bitwise.scala 48:55:@6143.4]
  wire [2:0] _T_6757; // @[Bitwise.scala 48:55:@6144.4]
  wire [3:0] _T_6758; // @[Bitwise.scala 48:55:@6145.4]
  wire [4:0] _T_6759; // @[Bitwise.scala 48:55:@6146.4]
  wire [5:0] _T_6760; // @[Bitwise.scala 48:55:@6147.4]
  wire [6:0] _T_6761; // @[Bitwise.scala 48:55:@6148.4]
  wire [50:0] _T_6825; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6213.4]
  wire  _T_6826; // @[Bitwise.scala 50:65:@6214.4]
  wire  _T_6827; // @[Bitwise.scala 50:65:@6215.4]
  wire  _T_6828; // @[Bitwise.scala 50:65:@6216.4]
  wire  _T_6829; // @[Bitwise.scala 50:65:@6217.4]
  wire  _T_6830; // @[Bitwise.scala 50:65:@6218.4]
  wire  _T_6831; // @[Bitwise.scala 50:65:@6219.4]
  wire  _T_6832; // @[Bitwise.scala 50:65:@6220.4]
  wire  _T_6833; // @[Bitwise.scala 50:65:@6221.4]
  wire  _T_6834; // @[Bitwise.scala 50:65:@6222.4]
  wire  _T_6835; // @[Bitwise.scala 50:65:@6223.4]
  wire  _T_6836; // @[Bitwise.scala 50:65:@6224.4]
  wire  _T_6837; // @[Bitwise.scala 50:65:@6225.4]
  wire  _T_6838; // @[Bitwise.scala 50:65:@6226.4]
  wire  _T_6839; // @[Bitwise.scala 50:65:@6227.4]
  wire  _T_6840; // @[Bitwise.scala 50:65:@6228.4]
  wire  _T_6841; // @[Bitwise.scala 50:65:@6229.4]
  wire  _T_6842; // @[Bitwise.scala 50:65:@6230.4]
  wire  _T_6843; // @[Bitwise.scala 50:65:@6231.4]
  wire  _T_6844; // @[Bitwise.scala 50:65:@6232.4]
  wire  _T_6845; // @[Bitwise.scala 50:65:@6233.4]
  wire  _T_6846; // @[Bitwise.scala 50:65:@6234.4]
  wire  _T_6847; // @[Bitwise.scala 50:65:@6235.4]
  wire  _T_6848; // @[Bitwise.scala 50:65:@6236.4]
  wire  _T_6849; // @[Bitwise.scala 50:65:@6237.4]
  wire  _T_6850; // @[Bitwise.scala 50:65:@6238.4]
  wire  _T_6851; // @[Bitwise.scala 50:65:@6239.4]
  wire  _T_6852; // @[Bitwise.scala 50:65:@6240.4]
  wire  _T_6853; // @[Bitwise.scala 50:65:@6241.4]
  wire  _T_6854; // @[Bitwise.scala 50:65:@6242.4]
  wire  _T_6855; // @[Bitwise.scala 50:65:@6243.4]
  wire  _T_6856; // @[Bitwise.scala 50:65:@6244.4]
  wire  _T_6857; // @[Bitwise.scala 50:65:@6245.4]
  wire  _T_6858; // @[Bitwise.scala 50:65:@6246.4]
  wire  _T_6859; // @[Bitwise.scala 50:65:@6247.4]
  wire  _T_6860; // @[Bitwise.scala 50:65:@6248.4]
  wire  _T_6861; // @[Bitwise.scala 50:65:@6249.4]
  wire  _T_6862; // @[Bitwise.scala 50:65:@6250.4]
  wire  _T_6863; // @[Bitwise.scala 50:65:@6251.4]
  wire  _T_6864; // @[Bitwise.scala 50:65:@6252.4]
  wire  _T_6865; // @[Bitwise.scala 50:65:@6253.4]
  wire  _T_6866; // @[Bitwise.scala 50:65:@6254.4]
  wire  _T_6867; // @[Bitwise.scala 50:65:@6255.4]
  wire  _T_6868; // @[Bitwise.scala 50:65:@6256.4]
  wire  _T_6869; // @[Bitwise.scala 50:65:@6257.4]
  wire  _T_6870; // @[Bitwise.scala 50:65:@6258.4]
  wire  _T_6871; // @[Bitwise.scala 50:65:@6259.4]
  wire  _T_6872; // @[Bitwise.scala 50:65:@6260.4]
  wire  _T_6873; // @[Bitwise.scala 50:65:@6261.4]
  wire  _T_6874; // @[Bitwise.scala 50:65:@6262.4]
  wire  _T_6875; // @[Bitwise.scala 50:65:@6263.4]
  wire  _T_6876; // @[Bitwise.scala 50:65:@6264.4]
  wire [1:0] _T_6877; // @[Bitwise.scala 48:55:@6265.4]
  wire [1:0] _GEN_906; // @[Bitwise.scala 48:55:@6266.4]
  wire [2:0] _T_6878; // @[Bitwise.scala 48:55:@6266.4]
  wire [1:0] _T_6879; // @[Bitwise.scala 48:55:@6267.4]
  wire [1:0] _GEN_907; // @[Bitwise.scala 48:55:@6268.4]
  wire [2:0] _T_6880; // @[Bitwise.scala 48:55:@6268.4]
  wire [3:0] _T_6881; // @[Bitwise.scala 48:55:@6269.4]
  wire [1:0] _T_6882; // @[Bitwise.scala 48:55:@6270.4]
  wire [1:0] _GEN_908; // @[Bitwise.scala 48:55:@6271.4]
  wire [2:0] _T_6883; // @[Bitwise.scala 48:55:@6271.4]
  wire [1:0] _T_6884; // @[Bitwise.scala 48:55:@6272.4]
  wire [1:0] _GEN_909; // @[Bitwise.scala 48:55:@6273.4]
  wire [2:0] _T_6885; // @[Bitwise.scala 48:55:@6273.4]
  wire [3:0] _T_6886; // @[Bitwise.scala 48:55:@6274.4]
  wire [4:0] _T_6887; // @[Bitwise.scala 48:55:@6275.4]
  wire [1:0] _T_6888; // @[Bitwise.scala 48:55:@6276.4]
  wire [1:0] _GEN_910; // @[Bitwise.scala 48:55:@6277.4]
  wire [2:0] _T_6889; // @[Bitwise.scala 48:55:@6277.4]
  wire [1:0] _T_6890; // @[Bitwise.scala 48:55:@6278.4]
  wire [1:0] _GEN_911; // @[Bitwise.scala 48:55:@6279.4]
  wire [2:0] _T_6891; // @[Bitwise.scala 48:55:@6279.4]
  wire [3:0] _T_6892; // @[Bitwise.scala 48:55:@6280.4]
  wire [1:0] _T_6893; // @[Bitwise.scala 48:55:@6281.4]
  wire [1:0] _GEN_912; // @[Bitwise.scala 48:55:@6282.4]
  wire [2:0] _T_6894; // @[Bitwise.scala 48:55:@6282.4]
  wire [1:0] _T_6895; // @[Bitwise.scala 48:55:@6283.4]
  wire [1:0] _T_6896; // @[Bitwise.scala 48:55:@6284.4]
  wire [2:0] _T_6897; // @[Bitwise.scala 48:55:@6285.4]
  wire [3:0] _T_6898; // @[Bitwise.scala 48:55:@6286.4]
  wire [4:0] _T_6899; // @[Bitwise.scala 48:55:@6287.4]
  wire [5:0] _T_6900; // @[Bitwise.scala 48:55:@6288.4]
  wire [1:0] _T_6901; // @[Bitwise.scala 48:55:@6289.4]
  wire [1:0] _GEN_913; // @[Bitwise.scala 48:55:@6290.4]
  wire [2:0] _T_6902; // @[Bitwise.scala 48:55:@6290.4]
  wire [1:0] _T_6903; // @[Bitwise.scala 48:55:@6291.4]
  wire [1:0] _GEN_914; // @[Bitwise.scala 48:55:@6292.4]
  wire [2:0] _T_6904; // @[Bitwise.scala 48:55:@6292.4]
  wire [3:0] _T_6905; // @[Bitwise.scala 48:55:@6293.4]
  wire [1:0] _T_6906; // @[Bitwise.scala 48:55:@6294.4]
  wire [1:0] _GEN_915; // @[Bitwise.scala 48:55:@6295.4]
  wire [2:0] _T_6907; // @[Bitwise.scala 48:55:@6295.4]
  wire [1:0] _T_6908; // @[Bitwise.scala 48:55:@6296.4]
  wire [1:0] _T_6909; // @[Bitwise.scala 48:55:@6297.4]
  wire [2:0] _T_6910; // @[Bitwise.scala 48:55:@6298.4]
  wire [3:0] _T_6911; // @[Bitwise.scala 48:55:@6299.4]
  wire [4:0] _T_6912; // @[Bitwise.scala 48:55:@6300.4]
  wire [1:0] _T_6913; // @[Bitwise.scala 48:55:@6301.4]
  wire [1:0] _GEN_916; // @[Bitwise.scala 48:55:@6302.4]
  wire [2:0] _T_6914; // @[Bitwise.scala 48:55:@6302.4]
  wire [1:0] _T_6915; // @[Bitwise.scala 48:55:@6303.4]
  wire [1:0] _GEN_917; // @[Bitwise.scala 48:55:@6304.4]
  wire [2:0] _T_6916; // @[Bitwise.scala 48:55:@6304.4]
  wire [3:0] _T_6917; // @[Bitwise.scala 48:55:@6305.4]
  wire [1:0] _T_6918; // @[Bitwise.scala 48:55:@6306.4]
  wire [1:0] _GEN_918; // @[Bitwise.scala 48:55:@6307.4]
  wire [2:0] _T_6919; // @[Bitwise.scala 48:55:@6307.4]
  wire [1:0] _T_6920; // @[Bitwise.scala 48:55:@6308.4]
  wire [1:0] _T_6921; // @[Bitwise.scala 48:55:@6309.4]
  wire [2:0] _T_6922; // @[Bitwise.scala 48:55:@6310.4]
  wire [3:0] _T_6923; // @[Bitwise.scala 48:55:@6311.4]
  wire [4:0] _T_6924; // @[Bitwise.scala 48:55:@6312.4]
  wire [5:0] _T_6925; // @[Bitwise.scala 48:55:@6313.4]
  wire [6:0] _T_6926; // @[Bitwise.scala 48:55:@6314.4]
  wire [51:0] _T_6990; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6379.4]
  wire  _T_6991; // @[Bitwise.scala 50:65:@6380.4]
  wire  _T_6992; // @[Bitwise.scala 50:65:@6381.4]
  wire  _T_6993; // @[Bitwise.scala 50:65:@6382.4]
  wire  _T_6994; // @[Bitwise.scala 50:65:@6383.4]
  wire  _T_6995; // @[Bitwise.scala 50:65:@6384.4]
  wire  _T_6996; // @[Bitwise.scala 50:65:@6385.4]
  wire  _T_6997; // @[Bitwise.scala 50:65:@6386.4]
  wire  _T_6998; // @[Bitwise.scala 50:65:@6387.4]
  wire  _T_6999; // @[Bitwise.scala 50:65:@6388.4]
  wire  _T_7000; // @[Bitwise.scala 50:65:@6389.4]
  wire  _T_7001; // @[Bitwise.scala 50:65:@6390.4]
  wire  _T_7002; // @[Bitwise.scala 50:65:@6391.4]
  wire  _T_7003; // @[Bitwise.scala 50:65:@6392.4]
  wire  _T_7004; // @[Bitwise.scala 50:65:@6393.4]
  wire  _T_7005; // @[Bitwise.scala 50:65:@6394.4]
  wire  _T_7006; // @[Bitwise.scala 50:65:@6395.4]
  wire  _T_7007; // @[Bitwise.scala 50:65:@6396.4]
  wire  _T_7008; // @[Bitwise.scala 50:65:@6397.4]
  wire  _T_7009; // @[Bitwise.scala 50:65:@6398.4]
  wire  _T_7010; // @[Bitwise.scala 50:65:@6399.4]
  wire  _T_7011; // @[Bitwise.scala 50:65:@6400.4]
  wire  _T_7012; // @[Bitwise.scala 50:65:@6401.4]
  wire  _T_7013; // @[Bitwise.scala 50:65:@6402.4]
  wire  _T_7014; // @[Bitwise.scala 50:65:@6403.4]
  wire  _T_7015; // @[Bitwise.scala 50:65:@6404.4]
  wire  _T_7016; // @[Bitwise.scala 50:65:@6405.4]
  wire  _T_7017; // @[Bitwise.scala 50:65:@6406.4]
  wire  _T_7018; // @[Bitwise.scala 50:65:@6407.4]
  wire  _T_7019; // @[Bitwise.scala 50:65:@6408.4]
  wire  _T_7020; // @[Bitwise.scala 50:65:@6409.4]
  wire  _T_7021; // @[Bitwise.scala 50:65:@6410.4]
  wire  _T_7022; // @[Bitwise.scala 50:65:@6411.4]
  wire  _T_7023; // @[Bitwise.scala 50:65:@6412.4]
  wire  _T_7024; // @[Bitwise.scala 50:65:@6413.4]
  wire  _T_7025; // @[Bitwise.scala 50:65:@6414.4]
  wire  _T_7026; // @[Bitwise.scala 50:65:@6415.4]
  wire  _T_7027; // @[Bitwise.scala 50:65:@6416.4]
  wire  _T_7028; // @[Bitwise.scala 50:65:@6417.4]
  wire  _T_7029; // @[Bitwise.scala 50:65:@6418.4]
  wire  _T_7030; // @[Bitwise.scala 50:65:@6419.4]
  wire  _T_7031; // @[Bitwise.scala 50:65:@6420.4]
  wire  _T_7032; // @[Bitwise.scala 50:65:@6421.4]
  wire  _T_7033; // @[Bitwise.scala 50:65:@6422.4]
  wire  _T_7034; // @[Bitwise.scala 50:65:@6423.4]
  wire  _T_7035; // @[Bitwise.scala 50:65:@6424.4]
  wire  _T_7036; // @[Bitwise.scala 50:65:@6425.4]
  wire  _T_7037; // @[Bitwise.scala 50:65:@6426.4]
  wire  _T_7038; // @[Bitwise.scala 50:65:@6427.4]
  wire  _T_7039; // @[Bitwise.scala 50:65:@6428.4]
  wire  _T_7040; // @[Bitwise.scala 50:65:@6429.4]
  wire  _T_7041; // @[Bitwise.scala 50:65:@6430.4]
  wire  _T_7042; // @[Bitwise.scala 50:65:@6431.4]
  wire [1:0] _T_7043; // @[Bitwise.scala 48:55:@6432.4]
  wire [1:0] _GEN_919; // @[Bitwise.scala 48:55:@6433.4]
  wire [2:0] _T_7044; // @[Bitwise.scala 48:55:@6433.4]
  wire [1:0] _T_7045; // @[Bitwise.scala 48:55:@6434.4]
  wire [1:0] _GEN_920; // @[Bitwise.scala 48:55:@6435.4]
  wire [2:0] _T_7046; // @[Bitwise.scala 48:55:@6435.4]
  wire [3:0] _T_7047; // @[Bitwise.scala 48:55:@6436.4]
  wire [1:0] _T_7048; // @[Bitwise.scala 48:55:@6437.4]
  wire [1:0] _GEN_921; // @[Bitwise.scala 48:55:@6438.4]
  wire [2:0] _T_7049; // @[Bitwise.scala 48:55:@6438.4]
  wire [1:0] _T_7050; // @[Bitwise.scala 48:55:@6439.4]
  wire [1:0] _T_7051; // @[Bitwise.scala 48:55:@6440.4]
  wire [2:0] _T_7052; // @[Bitwise.scala 48:55:@6441.4]
  wire [3:0] _T_7053; // @[Bitwise.scala 48:55:@6442.4]
  wire [4:0] _T_7054; // @[Bitwise.scala 48:55:@6443.4]
  wire [1:0] _T_7055; // @[Bitwise.scala 48:55:@6444.4]
  wire [1:0] _GEN_922; // @[Bitwise.scala 48:55:@6445.4]
  wire [2:0] _T_7056; // @[Bitwise.scala 48:55:@6445.4]
  wire [1:0] _T_7057; // @[Bitwise.scala 48:55:@6446.4]
  wire [1:0] _GEN_923; // @[Bitwise.scala 48:55:@6447.4]
  wire [2:0] _T_7058; // @[Bitwise.scala 48:55:@6447.4]
  wire [3:0] _T_7059; // @[Bitwise.scala 48:55:@6448.4]
  wire [1:0] _T_7060; // @[Bitwise.scala 48:55:@6449.4]
  wire [1:0] _GEN_924; // @[Bitwise.scala 48:55:@6450.4]
  wire [2:0] _T_7061; // @[Bitwise.scala 48:55:@6450.4]
  wire [1:0] _T_7062; // @[Bitwise.scala 48:55:@6451.4]
  wire [1:0] _T_7063; // @[Bitwise.scala 48:55:@6452.4]
  wire [2:0] _T_7064; // @[Bitwise.scala 48:55:@6453.4]
  wire [3:0] _T_7065; // @[Bitwise.scala 48:55:@6454.4]
  wire [4:0] _T_7066; // @[Bitwise.scala 48:55:@6455.4]
  wire [5:0] _T_7067; // @[Bitwise.scala 48:55:@6456.4]
  wire [1:0] _T_7068; // @[Bitwise.scala 48:55:@6457.4]
  wire [1:0] _GEN_925; // @[Bitwise.scala 48:55:@6458.4]
  wire [2:0] _T_7069; // @[Bitwise.scala 48:55:@6458.4]
  wire [1:0] _T_7070; // @[Bitwise.scala 48:55:@6459.4]
  wire [1:0] _GEN_926; // @[Bitwise.scala 48:55:@6460.4]
  wire [2:0] _T_7071; // @[Bitwise.scala 48:55:@6460.4]
  wire [3:0] _T_7072; // @[Bitwise.scala 48:55:@6461.4]
  wire [1:0] _T_7073; // @[Bitwise.scala 48:55:@6462.4]
  wire [1:0] _GEN_927; // @[Bitwise.scala 48:55:@6463.4]
  wire [2:0] _T_7074; // @[Bitwise.scala 48:55:@6463.4]
  wire [1:0] _T_7075; // @[Bitwise.scala 48:55:@6464.4]
  wire [1:0] _T_7076; // @[Bitwise.scala 48:55:@6465.4]
  wire [2:0] _T_7077; // @[Bitwise.scala 48:55:@6466.4]
  wire [3:0] _T_7078; // @[Bitwise.scala 48:55:@6467.4]
  wire [4:0] _T_7079; // @[Bitwise.scala 48:55:@6468.4]
  wire [1:0] _T_7080; // @[Bitwise.scala 48:55:@6469.4]
  wire [1:0] _GEN_928; // @[Bitwise.scala 48:55:@6470.4]
  wire [2:0] _T_7081; // @[Bitwise.scala 48:55:@6470.4]
  wire [1:0] _T_7082; // @[Bitwise.scala 48:55:@6471.4]
  wire [1:0] _GEN_929; // @[Bitwise.scala 48:55:@6472.4]
  wire [2:0] _T_7083; // @[Bitwise.scala 48:55:@6472.4]
  wire [3:0] _T_7084; // @[Bitwise.scala 48:55:@6473.4]
  wire [1:0] _T_7085; // @[Bitwise.scala 48:55:@6474.4]
  wire [1:0] _GEN_930; // @[Bitwise.scala 48:55:@6475.4]
  wire [2:0] _T_7086; // @[Bitwise.scala 48:55:@6475.4]
  wire [1:0] _T_7087; // @[Bitwise.scala 48:55:@6476.4]
  wire [1:0] _T_7088; // @[Bitwise.scala 48:55:@6477.4]
  wire [2:0] _T_7089; // @[Bitwise.scala 48:55:@6478.4]
  wire [3:0] _T_7090; // @[Bitwise.scala 48:55:@6479.4]
  wire [4:0] _T_7091; // @[Bitwise.scala 48:55:@6480.4]
  wire [5:0] _T_7092; // @[Bitwise.scala 48:55:@6481.4]
  wire [6:0] _T_7093; // @[Bitwise.scala 48:55:@6482.4]
  wire [52:0] _T_7157; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6547.4]
  wire  _T_7158; // @[Bitwise.scala 50:65:@6548.4]
  wire  _T_7159; // @[Bitwise.scala 50:65:@6549.4]
  wire  _T_7160; // @[Bitwise.scala 50:65:@6550.4]
  wire  _T_7161; // @[Bitwise.scala 50:65:@6551.4]
  wire  _T_7162; // @[Bitwise.scala 50:65:@6552.4]
  wire  _T_7163; // @[Bitwise.scala 50:65:@6553.4]
  wire  _T_7164; // @[Bitwise.scala 50:65:@6554.4]
  wire  _T_7165; // @[Bitwise.scala 50:65:@6555.4]
  wire  _T_7166; // @[Bitwise.scala 50:65:@6556.4]
  wire  _T_7167; // @[Bitwise.scala 50:65:@6557.4]
  wire  _T_7168; // @[Bitwise.scala 50:65:@6558.4]
  wire  _T_7169; // @[Bitwise.scala 50:65:@6559.4]
  wire  _T_7170; // @[Bitwise.scala 50:65:@6560.4]
  wire  _T_7171; // @[Bitwise.scala 50:65:@6561.4]
  wire  _T_7172; // @[Bitwise.scala 50:65:@6562.4]
  wire  _T_7173; // @[Bitwise.scala 50:65:@6563.4]
  wire  _T_7174; // @[Bitwise.scala 50:65:@6564.4]
  wire  _T_7175; // @[Bitwise.scala 50:65:@6565.4]
  wire  _T_7176; // @[Bitwise.scala 50:65:@6566.4]
  wire  _T_7177; // @[Bitwise.scala 50:65:@6567.4]
  wire  _T_7178; // @[Bitwise.scala 50:65:@6568.4]
  wire  _T_7179; // @[Bitwise.scala 50:65:@6569.4]
  wire  _T_7180; // @[Bitwise.scala 50:65:@6570.4]
  wire  _T_7181; // @[Bitwise.scala 50:65:@6571.4]
  wire  _T_7182; // @[Bitwise.scala 50:65:@6572.4]
  wire  _T_7183; // @[Bitwise.scala 50:65:@6573.4]
  wire  _T_7184; // @[Bitwise.scala 50:65:@6574.4]
  wire  _T_7185; // @[Bitwise.scala 50:65:@6575.4]
  wire  _T_7186; // @[Bitwise.scala 50:65:@6576.4]
  wire  _T_7187; // @[Bitwise.scala 50:65:@6577.4]
  wire  _T_7188; // @[Bitwise.scala 50:65:@6578.4]
  wire  _T_7189; // @[Bitwise.scala 50:65:@6579.4]
  wire  _T_7190; // @[Bitwise.scala 50:65:@6580.4]
  wire  _T_7191; // @[Bitwise.scala 50:65:@6581.4]
  wire  _T_7192; // @[Bitwise.scala 50:65:@6582.4]
  wire  _T_7193; // @[Bitwise.scala 50:65:@6583.4]
  wire  _T_7194; // @[Bitwise.scala 50:65:@6584.4]
  wire  _T_7195; // @[Bitwise.scala 50:65:@6585.4]
  wire  _T_7196; // @[Bitwise.scala 50:65:@6586.4]
  wire  _T_7197; // @[Bitwise.scala 50:65:@6587.4]
  wire  _T_7198; // @[Bitwise.scala 50:65:@6588.4]
  wire  _T_7199; // @[Bitwise.scala 50:65:@6589.4]
  wire  _T_7200; // @[Bitwise.scala 50:65:@6590.4]
  wire  _T_7201; // @[Bitwise.scala 50:65:@6591.4]
  wire  _T_7202; // @[Bitwise.scala 50:65:@6592.4]
  wire  _T_7203; // @[Bitwise.scala 50:65:@6593.4]
  wire  _T_7204; // @[Bitwise.scala 50:65:@6594.4]
  wire  _T_7205; // @[Bitwise.scala 50:65:@6595.4]
  wire  _T_7206; // @[Bitwise.scala 50:65:@6596.4]
  wire  _T_7207; // @[Bitwise.scala 50:65:@6597.4]
  wire  _T_7208; // @[Bitwise.scala 50:65:@6598.4]
  wire  _T_7209; // @[Bitwise.scala 50:65:@6599.4]
  wire  _T_7210; // @[Bitwise.scala 50:65:@6600.4]
  wire [1:0] _T_7211; // @[Bitwise.scala 48:55:@6601.4]
  wire [1:0] _GEN_931; // @[Bitwise.scala 48:55:@6602.4]
  wire [2:0] _T_7212; // @[Bitwise.scala 48:55:@6602.4]
  wire [1:0] _T_7213; // @[Bitwise.scala 48:55:@6603.4]
  wire [1:0] _GEN_932; // @[Bitwise.scala 48:55:@6604.4]
  wire [2:0] _T_7214; // @[Bitwise.scala 48:55:@6604.4]
  wire [3:0] _T_7215; // @[Bitwise.scala 48:55:@6605.4]
  wire [1:0] _T_7216; // @[Bitwise.scala 48:55:@6606.4]
  wire [1:0] _GEN_933; // @[Bitwise.scala 48:55:@6607.4]
  wire [2:0] _T_7217; // @[Bitwise.scala 48:55:@6607.4]
  wire [1:0] _T_7218; // @[Bitwise.scala 48:55:@6608.4]
  wire [1:0] _T_7219; // @[Bitwise.scala 48:55:@6609.4]
  wire [2:0] _T_7220; // @[Bitwise.scala 48:55:@6610.4]
  wire [3:0] _T_7221; // @[Bitwise.scala 48:55:@6611.4]
  wire [4:0] _T_7222; // @[Bitwise.scala 48:55:@6612.4]
  wire [1:0] _T_7223; // @[Bitwise.scala 48:55:@6613.4]
  wire [1:0] _GEN_934; // @[Bitwise.scala 48:55:@6614.4]
  wire [2:0] _T_7224; // @[Bitwise.scala 48:55:@6614.4]
  wire [1:0] _T_7225; // @[Bitwise.scala 48:55:@6615.4]
  wire [1:0] _GEN_935; // @[Bitwise.scala 48:55:@6616.4]
  wire [2:0] _T_7226; // @[Bitwise.scala 48:55:@6616.4]
  wire [3:0] _T_7227; // @[Bitwise.scala 48:55:@6617.4]
  wire [1:0] _T_7228; // @[Bitwise.scala 48:55:@6618.4]
  wire [1:0] _GEN_936; // @[Bitwise.scala 48:55:@6619.4]
  wire [2:0] _T_7229; // @[Bitwise.scala 48:55:@6619.4]
  wire [1:0] _T_7230; // @[Bitwise.scala 48:55:@6620.4]
  wire [1:0] _T_7231; // @[Bitwise.scala 48:55:@6621.4]
  wire [2:0] _T_7232; // @[Bitwise.scala 48:55:@6622.4]
  wire [3:0] _T_7233; // @[Bitwise.scala 48:55:@6623.4]
  wire [4:0] _T_7234; // @[Bitwise.scala 48:55:@6624.4]
  wire [5:0] _T_7235; // @[Bitwise.scala 48:55:@6625.4]
  wire [1:0] _T_7236; // @[Bitwise.scala 48:55:@6626.4]
  wire [1:0] _GEN_937; // @[Bitwise.scala 48:55:@6627.4]
  wire [2:0] _T_7237; // @[Bitwise.scala 48:55:@6627.4]
  wire [1:0] _T_7238; // @[Bitwise.scala 48:55:@6628.4]
  wire [1:0] _GEN_938; // @[Bitwise.scala 48:55:@6629.4]
  wire [2:0] _T_7239; // @[Bitwise.scala 48:55:@6629.4]
  wire [3:0] _T_7240; // @[Bitwise.scala 48:55:@6630.4]
  wire [1:0] _T_7241; // @[Bitwise.scala 48:55:@6631.4]
  wire [1:0] _GEN_939; // @[Bitwise.scala 48:55:@6632.4]
  wire [2:0] _T_7242; // @[Bitwise.scala 48:55:@6632.4]
  wire [1:0] _T_7243; // @[Bitwise.scala 48:55:@6633.4]
  wire [1:0] _T_7244; // @[Bitwise.scala 48:55:@6634.4]
  wire [2:0] _T_7245; // @[Bitwise.scala 48:55:@6635.4]
  wire [3:0] _T_7246; // @[Bitwise.scala 48:55:@6636.4]
  wire [4:0] _T_7247; // @[Bitwise.scala 48:55:@6637.4]
  wire [1:0] _T_7248; // @[Bitwise.scala 48:55:@6638.4]
  wire [1:0] _GEN_940; // @[Bitwise.scala 48:55:@6639.4]
  wire [2:0] _T_7249; // @[Bitwise.scala 48:55:@6639.4]
  wire [1:0] _T_7250; // @[Bitwise.scala 48:55:@6640.4]
  wire [1:0] _T_7251; // @[Bitwise.scala 48:55:@6641.4]
  wire [2:0] _T_7252; // @[Bitwise.scala 48:55:@6642.4]
  wire [3:0] _T_7253; // @[Bitwise.scala 48:55:@6643.4]
  wire [1:0] _T_7254; // @[Bitwise.scala 48:55:@6644.4]
  wire [1:0] _GEN_941; // @[Bitwise.scala 48:55:@6645.4]
  wire [2:0] _T_7255; // @[Bitwise.scala 48:55:@6645.4]
  wire [1:0] _T_7256; // @[Bitwise.scala 48:55:@6646.4]
  wire [1:0] _T_7257; // @[Bitwise.scala 48:55:@6647.4]
  wire [2:0] _T_7258; // @[Bitwise.scala 48:55:@6648.4]
  wire [3:0] _T_7259; // @[Bitwise.scala 48:55:@6649.4]
  wire [4:0] _T_7260; // @[Bitwise.scala 48:55:@6650.4]
  wire [5:0] _T_7261; // @[Bitwise.scala 48:55:@6651.4]
  wire [6:0] _T_7262; // @[Bitwise.scala 48:55:@6652.4]
  wire [53:0] _T_7326; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6717.4]
  wire  _T_7327; // @[Bitwise.scala 50:65:@6718.4]
  wire  _T_7328; // @[Bitwise.scala 50:65:@6719.4]
  wire  _T_7329; // @[Bitwise.scala 50:65:@6720.4]
  wire  _T_7330; // @[Bitwise.scala 50:65:@6721.4]
  wire  _T_7331; // @[Bitwise.scala 50:65:@6722.4]
  wire  _T_7332; // @[Bitwise.scala 50:65:@6723.4]
  wire  _T_7333; // @[Bitwise.scala 50:65:@6724.4]
  wire  _T_7334; // @[Bitwise.scala 50:65:@6725.4]
  wire  _T_7335; // @[Bitwise.scala 50:65:@6726.4]
  wire  _T_7336; // @[Bitwise.scala 50:65:@6727.4]
  wire  _T_7337; // @[Bitwise.scala 50:65:@6728.4]
  wire  _T_7338; // @[Bitwise.scala 50:65:@6729.4]
  wire  _T_7339; // @[Bitwise.scala 50:65:@6730.4]
  wire  _T_7340; // @[Bitwise.scala 50:65:@6731.4]
  wire  _T_7341; // @[Bitwise.scala 50:65:@6732.4]
  wire  _T_7342; // @[Bitwise.scala 50:65:@6733.4]
  wire  _T_7343; // @[Bitwise.scala 50:65:@6734.4]
  wire  _T_7344; // @[Bitwise.scala 50:65:@6735.4]
  wire  _T_7345; // @[Bitwise.scala 50:65:@6736.4]
  wire  _T_7346; // @[Bitwise.scala 50:65:@6737.4]
  wire  _T_7347; // @[Bitwise.scala 50:65:@6738.4]
  wire  _T_7348; // @[Bitwise.scala 50:65:@6739.4]
  wire  _T_7349; // @[Bitwise.scala 50:65:@6740.4]
  wire  _T_7350; // @[Bitwise.scala 50:65:@6741.4]
  wire  _T_7351; // @[Bitwise.scala 50:65:@6742.4]
  wire  _T_7352; // @[Bitwise.scala 50:65:@6743.4]
  wire  _T_7353; // @[Bitwise.scala 50:65:@6744.4]
  wire  _T_7354; // @[Bitwise.scala 50:65:@6745.4]
  wire  _T_7355; // @[Bitwise.scala 50:65:@6746.4]
  wire  _T_7356; // @[Bitwise.scala 50:65:@6747.4]
  wire  _T_7357; // @[Bitwise.scala 50:65:@6748.4]
  wire  _T_7358; // @[Bitwise.scala 50:65:@6749.4]
  wire  _T_7359; // @[Bitwise.scala 50:65:@6750.4]
  wire  _T_7360; // @[Bitwise.scala 50:65:@6751.4]
  wire  _T_7361; // @[Bitwise.scala 50:65:@6752.4]
  wire  _T_7362; // @[Bitwise.scala 50:65:@6753.4]
  wire  _T_7363; // @[Bitwise.scala 50:65:@6754.4]
  wire  _T_7364; // @[Bitwise.scala 50:65:@6755.4]
  wire  _T_7365; // @[Bitwise.scala 50:65:@6756.4]
  wire  _T_7366; // @[Bitwise.scala 50:65:@6757.4]
  wire  _T_7367; // @[Bitwise.scala 50:65:@6758.4]
  wire  _T_7368; // @[Bitwise.scala 50:65:@6759.4]
  wire  _T_7369; // @[Bitwise.scala 50:65:@6760.4]
  wire  _T_7370; // @[Bitwise.scala 50:65:@6761.4]
  wire  _T_7371; // @[Bitwise.scala 50:65:@6762.4]
  wire  _T_7372; // @[Bitwise.scala 50:65:@6763.4]
  wire  _T_7373; // @[Bitwise.scala 50:65:@6764.4]
  wire  _T_7374; // @[Bitwise.scala 50:65:@6765.4]
  wire  _T_7375; // @[Bitwise.scala 50:65:@6766.4]
  wire  _T_7376; // @[Bitwise.scala 50:65:@6767.4]
  wire  _T_7377; // @[Bitwise.scala 50:65:@6768.4]
  wire  _T_7378; // @[Bitwise.scala 50:65:@6769.4]
  wire  _T_7379; // @[Bitwise.scala 50:65:@6770.4]
  wire  _T_7380; // @[Bitwise.scala 50:65:@6771.4]
  wire [1:0] _T_7381; // @[Bitwise.scala 48:55:@6772.4]
  wire [1:0] _GEN_942; // @[Bitwise.scala 48:55:@6773.4]
  wire [2:0] _T_7382; // @[Bitwise.scala 48:55:@6773.4]
  wire [1:0] _T_7383; // @[Bitwise.scala 48:55:@6774.4]
  wire [1:0] _GEN_943; // @[Bitwise.scala 48:55:@6775.4]
  wire [2:0] _T_7384; // @[Bitwise.scala 48:55:@6775.4]
  wire [3:0] _T_7385; // @[Bitwise.scala 48:55:@6776.4]
  wire [1:0] _T_7386; // @[Bitwise.scala 48:55:@6777.4]
  wire [1:0] _GEN_944; // @[Bitwise.scala 48:55:@6778.4]
  wire [2:0] _T_7387; // @[Bitwise.scala 48:55:@6778.4]
  wire [1:0] _T_7388; // @[Bitwise.scala 48:55:@6779.4]
  wire [1:0] _T_7389; // @[Bitwise.scala 48:55:@6780.4]
  wire [2:0] _T_7390; // @[Bitwise.scala 48:55:@6781.4]
  wire [3:0] _T_7391; // @[Bitwise.scala 48:55:@6782.4]
  wire [4:0] _T_7392; // @[Bitwise.scala 48:55:@6783.4]
  wire [1:0] _T_7393; // @[Bitwise.scala 48:55:@6784.4]
  wire [1:0] _GEN_945; // @[Bitwise.scala 48:55:@6785.4]
  wire [2:0] _T_7394; // @[Bitwise.scala 48:55:@6785.4]
  wire [1:0] _T_7395; // @[Bitwise.scala 48:55:@6786.4]
  wire [1:0] _T_7396; // @[Bitwise.scala 48:55:@6787.4]
  wire [2:0] _T_7397; // @[Bitwise.scala 48:55:@6788.4]
  wire [3:0] _T_7398; // @[Bitwise.scala 48:55:@6789.4]
  wire [1:0] _T_7399; // @[Bitwise.scala 48:55:@6790.4]
  wire [1:0] _GEN_946; // @[Bitwise.scala 48:55:@6791.4]
  wire [2:0] _T_7400; // @[Bitwise.scala 48:55:@6791.4]
  wire [1:0] _T_7401; // @[Bitwise.scala 48:55:@6792.4]
  wire [1:0] _T_7402; // @[Bitwise.scala 48:55:@6793.4]
  wire [2:0] _T_7403; // @[Bitwise.scala 48:55:@6794.4]
  wire [3:0] _T_7404; // @[Bitwise.scala 48:55:@6795.4]
  wire [4:0] _T_7405; // @[Bitwise.scala 48:55:@6796.4]
  wire [5:0] _T_7406; // @[Bitwise.scala 48:55:@6797.4]
  wire [1:0] _T_7407; // @[Bitwise.scala 48:55:@6798.4]
  wire [1:0] _GEN_947; // @[Bitwise.scala 48:55:@6799.4]
  wire [2:0] _T_7408; // @[Bitwise.scala 48:55:@6799.4]
  wire [1:0] _T_7409; // @[Bitwise.scala 48:55:@6800.4]
  wire [1:0] _GEN_948; // @[Bitwise.scala 48:55:@6801.4]
  wire [2:0] _T_7410; // @[Bitwise.scala 48:55:@6801.4]
  wire [3:0] _T_7411; // @[Bitwise.scala 48:55:@6802.4]
  wire [1:0] _T_7412; // @[Bitwise.scala 48:55:@6803.4]
  wire [1:0] _GEN_949; // @[Bitwise.scala 48:55:@6804.4]
  wire [2:0] _T_7413; // @[Bitwise.scala 48:55:@6804.4]
  wire [1:0] _T_7414; // @[Bitwise.scala 48:55:@6805.4]
  wire [1:0] _T_7415; // @[Bitwise.scala 48:55:@6806.4]
  wire [2:0] _T_7416; // @[Bitwise.scala 48:55:@6807.4]
  wire [3:0] _T_7417; // @[Bitwise.scala 48:55:@6808.4]
  wire [4:0] _T_7418; // @[Bitwise.scala 48:55:@6809.4]
  wire [1:0] _T_7419; // @[Bitwise.scala 48:55:@6810.4]
  wire [1:0] _GEN_950; // @[Bitwise.scala 48:55:@6811.4]
  wire [2:0] _T_7420; // @[Bitwise.scala 48:55:@6811.4]
  wire [1:0] _T_7421; // @[Bitwise.scala 48:55:@6812.4]
  wire [1:0] _T_7422; // @[Bitwise.scala 48:55:@6813.4]
  wire [2:0] _T_7423; // @[Bitwise.scala 48:55:@6814.4]
  wire [3:0] _T_7424; // @[Bitwise.scala 48:55:@6815.4]
  wire [1:0] _T_7425; // @[Bitwise.scala 48:55:@6816.4]
  wire [1:0] _GEN_951; // @[Bitwise.scala 48:55:@6817.4]
  wire [2:0] _T_7426; // @[Bitwise.scala 48:55:@6817.4]
  wire [1:0] _T_7427; // @[Bitwise.scala 48:55:@6818.4]
  wire [1:0] _T_7428; // @[Bitwise.scala 48:55:@6819.4]
  wire [2:0] _T_7429; // @[Bitwise.scala 48:55:@6820.4]
  wire [3:0] _T_7430; // @[Bitwise.scala 48:55:@6821.4]
  wire [4:0] _T_7431; // @[Bitwise.scala 48:55:@6822.4]
  wire [5:0] _T_7432; // @[Bitwise.scala 48:55:@6823.4]
  wire [6:0] _T_7433; // @[Bitwise.scala 48:55:@6824.4]
  wire [54:0] _T_7497; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6889.4]
  wire  _T_7498; // @[Bitwise.scala 50:65:@6890.4]
  wire  _T_7499; // @[Bitwise.scala 50:65:@6891.4]
  wire  _T_7500; // @[Bitwise.scala 50:65:@6892.4]
  wire  _T_7501; // @[Bitwise.scala 50:65:@6893.4]
  wire  _T_7502; // @[Bitwise.scala 50:65:@6894.4]
  wire  _T_7503; // @[Bitwise.scala 50:65:@6895.4]
  wire  _T_7504; // @[Bitwise.scala 50:65:@6896.4]
  wire  _T_7505; // @[Bitwise.scala 50:65:@6897.4]
  wire  _T_7506; // @[Bitwise.scala 50:65:@6898.4]
  wire  _T_7507; // @[Bitwise.scala 50:65:@6899.4]
  wire  _T_7508; // @[Bitwise.scala 50:65:@6900.4]
  wire  _T_7509; // @[Bitwise.scala 50:65:@6901.4]
  wire  _T_7510; // @[Bitwise.scala 50:65:@6902.4]
  wire  _T_7511; // @[Bitwise.scala 50:65:@6903.4]
  wire  _T_7512; // @[Bitwise.scala 50:65:@6904.4]
  wire  _T_7513; // @[Bitwise.scala 50:65:@6905.4]
  wire  _T_7514; // @[Bitwise.scala 50:65:@6906.4]
  wire  _T_7515; // @[Bitwise.scala 50:65:@6907.4]
  wire  _T_7516; // @[Bitwise.scala 50:65:@6908.4]
  wire  _T_7517; // @[Bitwise.scala 50:65:@6909.4]
  wire  _T_7518; // @[Bitwise.scala 50:65:@6910.4]
  wire  _T_7519; // @[Bitwise.scala 50:65:@6911.4]
  wire  _T_7520; // @[Bitwise.scala 50:65:@6912.4]
  wire  _T_7521; // @[Bitwise.scala 50:65:@6913.4]
  wire  _T_7522; // @[Bitwise.scala 50:65:@6914.4]
  wire  _T_7523; // @[Bitwise.scala 50:65:@6915.4]
  wire  _T_7524; // @[Bitwise.scala 50:65:@6916.4]
  wire  _T_7525; // @[Bitwise.scala 50:65:@6917.4]
  wire  _T_7526; // @[Bitwise.scala 50:65:@6918.4]
  wire  _T_7527; // @[Bitwise.scala 50:65:@6919.4]
  wire  _T_7528; // @[Bitwise.scala 50:65:@6920.4]
  wire  _T_7529; // @[Bitwise.scala 50:65:@6921.4]
  wire  _T_7530; // @[Bitwise.scala 50:65:@6922.4]
  wire  _T_7531; // @[Bitwise.scala 50:65:@6923.4]
  wire  _T_7532; // @[Bitwise.scala 50:65:@6924.4]
  wire  _T_7533; // @[Bitwise.scala 50:65:@6925.4]
  wire  _T_7534; // @[Bitwise.scala 50:65:@6926.4]
  wire  _T_7535; // @[Bitwise.scala 50:65:@6927.4]
  wire  _T_7536; // @[Bitwise.scala 50:65:@6928.4]
  wire  _T_7537; // @[Bitwise.scala 50:65:@6929.4]
  wire  _T_7538; // @[Bitwise.scala 50:65:@6930.4]
  wire  _T_7539; // @[Bitwise.scala 50:65:@6931.4]
  wire  _T_7540; // @[Bitwise.scala 50:65:@6932.4]
  wire  _T_7541; // @[Bitwise.scala 50:65:@6933.4]
  wire  _T_7542; // @[Bitwise.scala 50:65:@6934.4]
  wire  _T_7543; // @[Bitwise.scala 50:65:@6935.4]
  wire  _T_7544; // @[Bitwise.scala 50:65:@6936.4]
  wire  _T_7545; // @[Bitwise.scala 50:65:@6937.4]
  wire  _T_7546; // @[Bitwise.scala 50:65:@6938.4]
  wire  _T_7547; // @[Bitwise.scala 50:65:@6939.4]
  wire  _T_7548; // @[Bitwise.scala 50:65:@6940.4]
  wire  _T_7549; // @[Bitwise.scala 50:65:@6941.4]
  wire  _T_7550; // @[Bitwise.scala 50:65:@6942.4]
  wire  _T_7551; // @[Bitwise.scala 50:65:@6943.4]
  wire  _T_7552; // @[Bitwise.scala 50:65:@6944.4]
  wire [1:0] _T_7553; // @[Bitwise.scala 48:55:@6945.4]
  wire [1:0] _GEN_952; // @[Bitwise.scala 48:55:@6946.4]
  wire [2:0] _T_7554; // @[Bitwise.scala 48:55:@6946.4]
  wire [1:0] _T_7555; // @[Bitwise.scala 48:55:@6947.4]
  wire [1:0] _GEN_953; // @[Bitwise.scala 48:55:@6948.4]
  wire [2:0] _T_7556; // @[Bitwise.scala 48:55:@6948.4]
  wire [3:0] _T_7557; // @[Bitwise.scala 48:55:@6949.4]
  wire [1:0] _T_7558; // @[Bitwise.scala 48:55:@6950.4]
  wire [1:0] _GEN_954; // @[Bitwise.scala 48:55:@6951.4]
  wire [2:0] _T_7559; // @[Bitwise.scala 48:55:@6951.4]
  wire [1:0] _T_7560; // @[Bitwise.scala 48:55:@6952.4]
  wire [1:0] _T_7561; // @[Bitwise.scala 48:55:@6953.4]
  wire [2:0] _T_7562; // @[Bitwise.scala 48:55:@6954.4]
  wire [3:0] _T_7563; // @[Bitwise.scala 48:55:@6955.4]
  wire [4:0] _T_7564; // @[Bitwise.scala 48:55:@6956.4]
  wire [1:0] _T_7565; // @[Bitwise.scala 48:55:@6957.4]
  wire [1:0] _GEN_955; // @[Bitwise.scala 48:55:@6958.4]
  wire [2:0] _T_7566; // @[Bitwise.scala 48:55:@6958.4]
  wire [1:0] _T_7567; // @[Bitwise.scala 48:55:@6959.4]
  wire [1:0] _T_7568; // @[Bitwise.scala 48:55:@6960.4]
  wire [2:0] _T_7569; // @[Bitwise.scala 48:55:@6961.4]
  wire [3:0] _T_7570; // @[Bitwise.scala 48:55:@6962.4]
  wire [1:0] _T_7571; // @[Bitwise.scala 48:55:@6963.4]
  wire [1:0] _GEN_956; // @[Bitwise.scala 48:55:@6964.4]
  wire [2:0] _T_7572; // @[Bitwise.scala 48:55:@6964.4]
  wire [1:0] _T_7573; // @[Bitwise.scala 48:55:@6965.4]
  wire [1:0] _T_7574; // @[Bitwise.scala 48:55:@6966.4]
  wire [2:0] _T_7575; // @[Bitwise.scala 48:55:@6967.4]
  wire [3:0] _T_7576; // @[Bitwise.scala 48:55:@6968.4]
  wire [4:0] _T_7577; // @[Bitwise.scala 48:55:@6969.4]
  wire [5:0] _T_7578; // @[Bitwise.scala 48:55:@6970.4]
  wire [1:0] _T_7579; // @[Bitwise.scala 48:55:@6971.4]
  wire [1:0] _GEN_957; // @[Bitwise.scala 48:55:@6972.4]
  wire [2:0] _T_7580; // @[Bitwise.scala 48:55:@6972.4]
  wire [1:0] _T_7581; // @[Bitwise.scala 48:55:@6973.4]
  wire [1:0] _T_7582; // @[Bitwise.scala 48:55:@6974.4]
  wire [2:0] _T_7583; // @[Bitwise.scala 48:55:@6975.4]
  wire [3:0] _T_7584; // @[Bitwise.scala 48:55:@6976.4]
  wire [1:0] _T_7585; // @[Bitwise.scala 48:55:@6977.4]
  wire [1:0] _GEN_958; // @[Bitwise.scala 48:55:@6978.4]
  wire [2:0] _T_7586; // @[Bitwise.scala 48:55:@6978.4]
  wire [1:0] _T_7587; // @[Bitwise.scala 48:55:@6979.4]
  wire [1:0] _T_7588; // @[Bitwise.scala 48:55:@6980.4]
  wire [2:0] _T_7589; // @[Bitwise.scala 48:55:@6981.4]
  wire [3:0] _T_7590; // @[Bitwise.scala 48:55:@6982.4]
  wire [4:0] _T_7591; // @[Bitwise.scala 48:55:@6983.4]
  wire [1:0] _T_7592; // @[Bitwise.scala 48:55:@6984.4]
  wire [1:0] _GEN_959; // @[Bitwise.scala 48:55:@6985.4]
  wire [2:0] _T_7593; // @[Bitwise.scala 48:55:@6985.4]
  wire [1:0] _T_7594; // @[Bitwise.scala 48:55:@6986.4]
  wire [1:0] _T_7595; // @[Bitwise.scala 48:55:@6987.4]
  wire [2:0] _T_7596; // @[Bitwise.scala 48:55:@6988.4]
  wire [3:0] _T_7597; // @[Bitwise.scala 48:55:@6989.4]
  wire [1:0] _T_7598; // @[Bitwise.scala 48:55:@6990.4]
  wire [1:0] _GEN_960; // @[Bitwise.scala 48:55:@6991.4]
  wire [2:0] _T_7599; // @[Bitwise.scala 48:55:@6991.4]
  wire [1:0] _T_7600; // @[Bitwise.scala 48:55:@6992.4]
  wire [1:0] _T_7601; // @[Bitwise.scala 48:55:@6993.4]
  wire [2:0] _T_7602; // @[Bitwise.scala 48:55:@6994.4]
  wire [3:0] _T_7603; // @[Bitwise.scala 48:55:@6995.4]
  wire [4:0] _T_7604; // @[Bitwise.scala 48:55:@6996.4]
  wire [5:0] _T_7605; // @[Bitwise.scala 48:55:@6997.4]
  wire [6:0] _T_7606; // @[Bitwise.scala 48:55:@6998.4]
  wire [55:0] _T_7670; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7063.4]
  wire  _T_7671; // @[Bitwise.scala 50:65:@7064.4]
  wire  _T_7672; // @[Bitwise.scala 50:65:@7065.4]
  wire  _T_7673; // @[Bitwise.scala 50:65:@7066.4]
  wire  _T_7674; // @[Bitwise.scala 50:65:@7067.4]
  wire  _T_7675; // @[Bitwise.scala 50:65:@7068.4]
  wire  _T_7676; // @[Bitwise.scala 50:65:@7069.4]
  wire  _T_7677; // @[Bitwise.scala 50:65:@7070.4]
  wire  _T_7678; // @[Bitwise.scala 50:65:@7071.4]
  wire  _T_7679; // @[Bitwise.scala 50:65:@7072.4]
  wire  _T_7680; // @[Bitwise.scala 50:65:@7073.4]
  wire  _T_7681; // @[Bitwise.scala 50:65:@7074.4]
  wire  _T_7682; // @[Bitwise.scala 50:65:@7075.4]
  wire  _T_7683; // @[Bitwise.scala 50:65:@7076.4]
  wire  _T_7684; // @[Bitwise.scala 50:65:@7077.4]
  wire  _T_7685; // @[Bitwise.scala 50:65:@7078.4]
  wire  _T_7686; // @[Bitwise.scala 50:65:@7079.4]
  wire  _T_7687; // @[Bitwise.scala 50:65:@7080.4]
  wire  _T_7688; // @[Bitwise.scala 50:65:@7081.4]
  wire  _T_7689; // @[Bitwise.scala 50:65:@7082.4]
  wire  _T_7690; // @[Bitwise.scala 50:65:@7083.4]
  wire  _T_7691; // @[Bitwise.scala 50:65:@7084.4]
  wire  _T_7692; // @[Bitwise.scala 50:65:@7085.4]
  wire  _T_7693; // @[Bitwise.scala 50:65:@7086.4]
  wire  _T_7694; // @[Bitwise.scala 50:65:@7087.4]
  wire  _T_7695; // @[Bitwise.scala 50:65:@7088.4]
  wire  _T_7696; // @[Bitwise.scala 50:65:@7089.4]
  wire  _T_7697; // @[Bitwise.scala 50:65:@7090.4]
  wire  _T_7698; // @[Bitwise.scala 50:65:@7091.4]
  wire  _T_7699; // @[Bitwise.scala 50:65:@7092.4]
  wire  _T_7700; // @[Bitwise.scala 50:65:@7093.4]
  wire  _T_7701; // @[Bitwise.scala 50:65:@7094.4]
  wire  _T_7702; // @[Bitwise.scala 50:65:@7095.4]
  wire  _T_7703; // @[Bitwise.scala 50:65:@7096.4]
  wire  _T_7704; // @[Bitwise.scala 50:65:@7097.4]
  wire  _T_7705; // @[Bitwise.scala 50:65:@7098.4]
  wire  _T_7706; // @[Bitwise.scala 50:65:@7099.4]
  wire  _T_7707; // @[Bitwise.scala 50:65:@7100.4]
  wire  _T_7708; // @[Bitwise.scala 50:65:@7101.4]
  wire  _T_7709; // @[Bitwise.scala 50:65:@7102.4]
  wire  _T_7710; // @[Bitwise.scala 50:65:@7103.4]
  wire  _T_7711; // @[Bitwise.scala 50:65:@7104.4]
  wire  _T_7712; // @[Bitwise.scala 50:65:@7105.4]
  wire  _T_7713; // @[Bitwise.scala 50:65:@7106.4]
  wire  _T_7714; // @[Bitwise.scala 50:65:@7107.4]
  wire  _T_7715; // @[Bitwise.scala 50:65:@7108.4]
  wire  _T_7716; // @[Bitwise.scala 50:65:@7109.4]
  wire  _T_7717; // @[Bitwise.scala 50:65:@7110.4]
  wire  _T_7718; // @[Bitwise.scala 50:65:@7111.4]
  wire  _T_7719; // @[Bitwise.scala 50:65:@7112.4]
  wire  _T_7720; // @[Bitwise.scala 50:65:@7113.4]
  wire  _T_7721; // @[Bitwise.scala 50:65:@7114.4]
  wire  _T_7722; // @[Bitwise.scala 50:65:@7115.4]
  wire  _T_7723; // @[Bitwise.scala 50:65:@7116.4]
  wire  _T_7724; // @[Bitwise.scala 50:65:@7117.4]
  wire  _T_7725; // @[Bitwise.scala 50:65:@7118.4]
  wire  _T_7726; // @[Bitwise.scala 50:65:@7119.4]
  wire [1:0] _T_7727; // @[Bitwise.scala 48:55:@7120.4]
  wire [1:0] _GEN_961; // @[Bitwise.scala 48:55:@7121.4]
  wire [2:0] _T_7728; // @[Bitwise.scala 48:55:@7121.4]
  wire [1:0] _T_7729; // @[Bitwise.scala 48:55:@7122.4]
  wire [1:0] _T_7730; // @[Bitwise.scala 48:55:@7123.4]
  wire [2:0] _T_7731; // @[Bitwise.scala 48:55:@7124.4]
  wire [3:0] _T_7732; // @[Bitwise.scala 48:55:@7125.4]
  wire [1:0] _T_7733; // @[Bitwise.scala 48:55:@7126.4]
  wire [1:0] _GEN_962; // @[Bitwise.scala 48:55:@7127.4]
  wire [2:0] _T_7734; // @[Bitwise.scala 48:55:@7127.4]
  wire [1:0] _T_7735; // @[Bitwise.scala 48:55:@7128.4]
  wire [1:0] _T_7736; // @[Bitwise.scala 48:55:@7129.4]
  wire [2:0] _T_7737; // @[Bitwise.scala 48:55:@7130.4]
  wire [3:0] _T_7738; // @[Bitwise.scala 48:55:@7131.4]
  wire [4:0] _T_7739; // @[Bitwise.scala 48:55:@7132.4]
  wire [1:0] _T_7740; // @[Bitwise.scala 48:55:@7133.4]
  wire [1:0] _GEN_963; // @[Bitwise.scala 48:55:@7134.4]
  wire [2:0] _T_7741; // @[Bitwise.scala 48:55:@7134.4]
  wire [1:0] _T_7742; // @[Bitwise.scala 48:55:@7135.4]
  wire [1:0] _T_7743; // @[Bitwise.scala 48:55:@7136.4]
  wire [2:0] _T_7744; // @[Bitwise.scala 48:55:@7137.4]
  wire [3:0] _T_7745; // @[Bitwise.scala 48:55:@7138.4]
  wire [1:0] _T_7746; // @[Bitwise.scala 48:55:@7139.4]
  wire [1:0] _GEN_964; // @[Bitwise.scala 48:55:@7140.4]
  wire [2:0] _T_7747; // @[Bitwise.scala 48:55:@7140.4]
  wire [1:0] _T_7748; // @[Bitwise.scala 48:55:@7141.4]
  wire [1:0] _T_7749; // @[Bitwise.scala 48:55:@7142.4]
  wire [2:0] _T_7750; // @[Bitwise.scala 48:55:@7143.4]
  wire [3:0] _T_7751; // @[Bitwise.scala 48:55:@7144.4]
  wire [4:0] _T_7752; // @[Bitwise.scala 48:55:@7145.4]
  wire [5:0] _T_7753; // @[Bitwise.scala 48:55:@7146.4]
  wire [1:0] _T_7754; // @[Bitwise.scala 48:55:@7147.4]
  wire [1:0] _GEN_965; // @[Bitwise.scala 48:55:@7148.4]
  wire [2:0] _T_7755; // @[Bitwise.scala 48:55:@7148.4]
  wire [1:0] _T_7756; // @[Bitwise.scala 48:55:@7149.4]
  wire [1:0] _T_7757; // @[Bitwise.scala 48:55:@7150.4]
  wire [2:0] _T_7758; // @[Bitwise.scala 48:55:@7151.4]
  wire [3:0] _T_7759; // @[Bitwise.scala 48:55:@7152.4]
  wire [1:0] _T_7760; // @[Bitwise.scala 48:55:@7153.4]
  wire [1:0] _GEN_966; // @[Bitwise.scala 48:55:@7154.4]
  wire [2:0] _T_7761; // @[Bitwise.scala 48:55:@7154.4]
  wire [1:0] _T_7762; // @[Bitwise.scala 48:55:@7155.4]
  wire [1:0] _T_7763; // @[Bitwise.scala 48:55:@7156.4]
  wire [2:0] _T_7764; // @[Bitwise.scala 48:55:@7157.4]
  wire [3:0] _T_7765; // @[Bitwise.scala 48:55:@7158.4]
  wire [4:0] _T_7766; // @[Bitwise.scala 48:55:@7159.4]
  wire [1:0] _T_7767; // @[Bitwise.scala 48:55:@7160.4]
  wire [1:0] _GEN_967; // @[Bitwise.scala 48:55:@7161.4]
  wire [2:0] _T_7768; // @[Bitwise.scala 48:55:@7161.4]
  wire [1:0] _T_7769; // @[Bitwise.scala 48:55:@7162.4]
  wire [1:0] _T_7770; // @[Bitwise.scala 48:55:@7163.4]
  wire [2:0] _T_7771; // @[Bitwise.scala 48:55:@7164.4]
  wire [3:0] _T_7772; // @[Bitwise.scala 48:55:@7165.4]
  wire [1:0] _T_7773; // @[Bitwise.scala 48:55:@7166.4]
  wire [1:0] _GEN_968; // @[Bitwise.scala 48:55:@7167.4]
  wire [2:0] _T_7774; // @[Bitwise.scala 48:55:@7167.4]
  wire [1:0] _T_7775; // @[Bitwise.scala 48:55:@7168.4]
  wire [1:0] _T_7776; // @[Bitwise.scala 48:55:@7169.4]
  wire [2:0] _T_7777; // @[Bitwise.scala 48:55:@7170.4]
  wire [3:0] _T_7778; // @[Bitwise.scala 48:55:@7171.4]
  wire [4:0] _T_7779; // @[Bitwise.scala 48:55:@7172.4]
  wire [5:0] _T_7780; // @[Bitwise.scala 48:55:@7173.4]
  wire [6:0] _T_7781; // @[Bitwise.scala 48:55:@7174.4]
  wire [56:0] _T_7845; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7239.4]
  wire  _T_7846; // @[Bitwise.scala 50:65:@7240.4]
  wire  _T_7847; // @[Bitwise.scala 50:65:@7241.4]
  wire  _T_7848; // @[Bitwise.scala 50:65:@7242.4]
  wire  _T_7849; // @[Bitwise.scala 50:65:@7243.4]
  wire  _T_7850; // @[Bitwise.scala 50:65:@7244.4]
  wire  _T_7851; // @[Bitwise.scala 50:65:@7245.4]
  wire  _T_7852; // @[Bitwise.scala 50:65:@7246.4]
  wire  _T_7853; // @[Bitwise.scala 50:65:@7247.4]
  wire  _T_7854; // @[Bitwise.scala 50:65:@7248.4]
  wire  _T_7855; // @[Bitwise.scala 50:65:@7249.4]
  wire  _T_7856; // @[Bitwise.scala 50:65:@7250.4]
  wire  _T_7857; // @[Bitwise.scala 50:65:@7251.4]
  wire  _T_7858; // @[Bitwise.scala 50:65:@7252.4]
  wire  _T_7859; // @[Bitwise.scala 50:65:@7253.4]
  wire  _T_7860; // @[Bitwise.scala 50:65:@7254.4]
  wire  _T_7861; // @[Bitwise.scala 50:65:@7255.4]
  wire  _T_7862; // @[Bitwise.scala 50:65:@7256.4]
  wire  _T_7863; // @[Bitwise.scala 50:65:@7257.4]
  wire  _T_7864; // @[Bitwise.scala 50:65:@7258.4]
  wire  _T_7865; // @[Bitwise.scala 50:65:@7259.4]
  wire  _T_7866; // @[Bitwise.scala 50:65:@7260.4]
  wire  _T_7867; // @[Bitwise.scala 50:65:@7261.4]
  wire  _T_7868; // @[Bitwise.scala 50:65:@7262.4]
  wire  _T_7869; // @[Bitwise.scala 50:65:@7263.4]
  wire  _T_7870; // @[Bitwise.scala 50:65:@7264.4]
  wire  _T_7871; // @[Bitwise.scala 50:65:@7265.4]
  wire  _T_7872; // @[Bitwise.scala 50:65:@7266.4]
  wire  _T_7873; // @[Bitwise.scala 50:65:@7267.4]
  wire  _T_7874; // @[Bitwise.scala 50:65:@7268.4]
  wire  _T_7875; // @[Bitwise.scala 50:65:@7269.4]
  wire  _T_7876; // @[Bitwise.scala 50:65:@7270.4]
  wire  _T_7877; // @[Bitwise.scala 50:65:@7271.4]
  wire  _T_7878; // @[Bitwise.scala 50:65:@7272.4]
  wire  _T_7879; // @[Bitwise.scala 50:65:@7273.4]
  wire  _T_7880; // @[Bitwise.scala 50:65:@7274.4]
  wire  _T_7881; // @[Bitwise.scala 50:65:@7275.4]
  wire  _T_7882; // @[Bitwise.scala 50:65:@7276.4]
  wire  _T_7883; // @[Bitwise.scala 50:65:@7277.4]
  wire  _T_7884; // @[Bitwise.scala 50:65:@7278.4]
  wire  _T_7885; // @[Bitwise.scala 50:65:@7279.4]
  wire  _T_7886; // @[Bitwise.scala 50:65:@7280.4]
  wire  _T_7887; // @[Bitwise.scala 50:65:@7281.4]
  wire  _T_7888; // @[Bitwise.scala 50:65:@7282.4]
  wire  _T_7889; // @[Bitwise.scala 50:65:@7283.4]
  wire  _T_7890; // @[Bitwise.scala 50:65:@7284.4]
  wire  _T_7891; // @[Bitwise.scala 50:65:@7285.4]
  wire  _T_7892; // @[Bitwise.scala 50:65:@7286.4]
  wire  _T_7893; // @[Bitwise.scala 50:65:@7287.4]
  wire  _T_7894; // @[Bitwise.scala 50:65:@7288.4]
  wire  _T_7895; // @[Bitwise.scala 50:65:@7289.4]
  wire  _T_7896; // @[Bitwise.scala 50:65:@7290.4]
  wire  _T_7897; // @[Bitwise.scala 50:65:@7291.4]
  wire  _T_7898; // @[Bitwise.scala 50:65:@7292.4]
  wire  _T_7899; // @[Bitwise.scala 50:65:@7293.4]
  wire  _T_7900; // @[Bitwise.scala 50:65:@7294.4]
  wire  _T_7901; // @[Bitwise.scala 50:65:@7295.4]
  wire  _T_7902; // @[Bitwise.scala 50:65:@7296.4]
  wire [1:0] _T_7903; // @[Bitwise.scala 48:55:@7297.4]
  wire [1:0] _GEN_969; // @[Bitwise.scala 48:55:@7298.4]
  wire [2:0] _T_7904; // @[Bitwise.scala 48:55:@7298.4]
  wire [1:0] _T_7905; // @[Bitwise.scala 48:55:@7299.4]
  wire [1:0] _T_7906; // @[Bitwise.scala 48:55:@7300.4]
  wire [2:0] _T_7907; // @[Bitwise.scala 48:55:@7301.4]
  wire [3:0] _T_7908; // @[Bitwise.scala 48:55:@7302.4]
  wire [1:0] _T_7909; // @[Bitwise.scala 48:55:@7303.4]
  wire [1:0] _GEN_970; // @[Bitwise.scala 48:55:@7304.4]
  wire [2:0] _T_7910; // @[Bitwise.scala 48:55:@7304.4]
  wire [1:0] _T_7911; // @[Bitwise.scala 48:55:@7305.4]
  wire [1:0] _T_7912; // @[Bitwise.scala 48:55:@7306.4]
  wire [2:0] _T_7913; // @[Bitwise.scala 48:55:@7307.4]
  wire [3:0] _T_7914; // @[Bitwise.scala 48:55:@7308.4]
  wire [4:0] _T_7915; // @[Bitwise.scala 48:55:@7309.4]
  wire [1:0] _T_7916; // @[Bitwise.scala 48:55:@7310.4]
  wire [1:0] _GEN_971; // @[Bitwise.scala 48:55:@7311.4]
  wire [2:0] _T_7917; // @[Bitwise.scala 48:55:@7311.4]
  wire [1:0] _T_7918; // @[Bitwise.scala 48:55:@7312.4]
  wire [1:0] _T_7919; // @[Bitwise.scala 48:55:@7313.4]
  wire [2:0] _T_7920; // @[Bitwise.scala 48:55:@7314.4]
  wire [3:0] _T_7921; // @[Bitwise.scala 48:55:@7315.4]
  wire [1:0] _T_7922; // @[Bitwise.scala 48:55:@7316.4]
  wire [1:0] _GEN_972; // @[Bitwise.scala 48:55:@7317.4]
  wire [2:0] _T_7923; // @[Bitwise.scala 48:55:@7317.4]
  wire [1:0] _T_7924; // @[Bitwise.scala 48:55:@7318.4]
  wire [1:0] _T_7925; // @[Bitwise.scala 48:55:@7319.4]
  wire [2:0] _T_7926; // @[Bitwise.scala 48:55:@7320.4]
  wire [3:0] _T_7927; // @[Bitwise.scala 48:55:@7321.4]
  wire [4:0] _T_7928; // @[Bitwise.scala 48:55:@7322.4]
  wire [5:0] _T_7929; // @[Bitwise.scala 48:55:@7323.4]
  wire [1:0] _T_7930; // @[Bitwise.scala 48:55:@7324.4]
  wire [1:0] _GEN_973; // @[Bitwise.scala 48:55:@7325.4]
  wire [2:0] _T_7931; // @[Bitwise.scala 48:55:@7325.4]
  wire [1:0] _T_7932; // @[Bitwise.scala 48:55:@7326.4]
  wire [1:0] _T_7933; // @[Bitwise.scala 48:55:@7327.4]
  wire [2:0] _T_7934; // @[Bitwise.scala 48:55:@7328.4]
  wire [3:0] _T_7935; // @[Bitwise.scala 48:55:@7329.4]
  wire [1:0] _T_7936; // @[Bitwise.scala 48:55:@7330.4]
  wire [1:0] _GEN_974; // @[Bitwise.scala 48:55:@7331.4]
  wire [2:0] _T_7937; // @[Bitwise.scala 48:55:@7331.4]
  wire [1:0] _T_7938; // @[Bitwise.scala 48:55:@7332.4]
  wire [1:0] _T_7939; // @[Bitwise.scala 48:55:@7333.4]
  wire [2:0] _T_7940; // @[Bitwise.scala 48:55:@7334.4]
  wire [3:0] _T_7941; // @[Bitwise.scala 48:55:@7335.4]
  wire [4:0] _T_7942; // @[Bitwise.scala 48:55:@7336.4]
  wire [1:0] _T_7943; // @[Bitwise.scala 48:55:@7337.4]
  wire [1:0] _GEN_975; // @[Bitwise.scala 48:55:@7338.4]
  wire [2:0] _T_7944; // @[Bitwise.scala 48:55:@7338.4]
  wire [1:0] _T_7945; // @[Bitwise.scala 48:55:@7339.4]
  wire [1:0] _T_7946; // @[Bitwise.scala 48:55:@7340.4]
  wire [2:0] _T_7947; // @[Bitwise.scala 48:55:@7341.4]
  wire [3:0] _T_7948; // @[Bitwise.scala 48:55:@7342.4]
  wire [1:0] _T_7949; // @[Bitwise.scala 48:55:@7343.4]
  wire [1:0] _T_7950; // @[Bitwise.scala 48:55:@7344.4]
  wire [2:0] _T_7951; // @[Bitwise.scala 48:55:@7345.4]
  wire [1:0] _T_7952; // @[Bitwise.scala 48:55:@7346.4]
  wire [1:0] _T_7953; // @[Bitwise.scala 48:55:@7347.4]
  wire [2:0] _T_7954; // @[Bitwise.scala 48:55:@7348.4]
  wire [3:0] _T_7955; // @[Bitwise.scala 48:55:@7349.4]
  wire [4:0] _T_7956; // @[Bitwise.scala 48:55:@7350.4]
  wire [5:0] _T_7957; // @[Bitwise.scala 48:55:@7351.4]
  wire [6:0] _T_7958; // @[Bitwise.scala 48:55:@7352.4]
  wire [57:0] _T_8022; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7417.4]
  wire  _T_8023; // @[Bitwise.scala 50:65:@7418.4]
  wire  _T_8024; // @[Bitwise.scala 50:65:@7419.4]
  wire  _T_8025; // @[Bitwise.scala 50:65:@7420.4]
  wire  _T_8026; // @[Bitwise.scala 50:65:@7421.4]
  wire  _T_8027; // @[Bitwise.scala 50:65:@7422.4]
  wire  _T_8028; // @[Bitwise.scala 50:65:@7423.4]
  wire  _T_8029; // @[Bitwise.scala 50:65:@7424.4]
  wire  _T_8030; // @[Bitwise.scala 50:65:@7425.4]
  wire  _T_8031; // @[Bitwise.scala 50:65:@7426.4]
  wire  _T_8032; // @[Bitwise.scala 50:65:@7427.4]
  wire  _T_8033; // @[Bitwise.scala 50:65:@7428.4]
  wire  _T_8034; // @[Bitwise.scala 50:65:@7429.4]
  wire  _T_8035; // @[Bitwise.scala 50:65:@7430.4]
  wire  _T_8036; // @[Bitwise.scala 50:65:@7431.4]
  wire  _T_8037; // @[Bitwise.scala 50:65:@7432.4]
  wire  _T_8038; // @[Bitwise.scala 50:65:@7433.4]
  wire  _T_8039; // @[Bitwise.scala 50:65:@7434.4]
  wire  _T_8040; // @[Bitwise.scala 50:65:@7435.4]
  wire  _T_8041; // @[Bitwise.scala 50:65:@7436.4]
  wire  _T_8042; // @[Bitwise.scala 50:65:@7437.4]
  wire  _T_8043; // @[Bitwise.scala 50:65:@7438.4]
  wire  _T_8044; // @[Bitwise.scala 50:65:@7439.4]
  wire  _T_8045; // @[Bitwise.scala 50:65:@7440.4]
  wire  _T_8046; // @[Bitwise.scala 50:65:@7441.4]
  wire  _T_8047; // @[Bitwise.scala 50:65:@7442.4]
  wire  _T_8048; // @[Bitwise.scala 50:65:@7443.4]
  wire  _T_8049; // @[Bitwise.scala 50:65:@7444.4]
  wire  _T_8050; // @[Bitwise.scala 50:65:@7445.4]
  wire  _T_8051; // @[Bitwise.scala 50:65:@7446.4]
  wire  _T_8052; // @[Bitwise.scala 50:65:@7447.4]
  wire  _T_8053; // @[Bitwise.scala 50:65:@7448.4]
  wire  _T_8054; // @[Bitwise.scala 50:65:@7449.4]
  wire  _T_8055; // @[Bitwise.scala 50:65:@7450.4]
  wire  _T_8056; // @[Bitwise.scala 50:65:@7451.4]
  wire  _T_8057; // @[Bitwise.scala 50:65:@7452.4]
  wire  _T_8058; // @[Bitwise.scala 50:65:@7453.4]
  wire  _T_8059; // @[Bitwise.scala 50:65:@7454.4]
  wire  _T_8060; // @[Bitwise.scala 50:65:@7455.4]
  wire  _T_8061; // @[Bitwise.scala 50:65:@7456.4]
  wire  _T_8062; // @[Bitwise.scala 50:65:@7457.4]
  wire  _T_8063; // @[Bitwise.scala 50:65:@7458.4]
  wire  _T_8064; // @[Bitwise.scala 50:65:@7459.4]
  wire  _T_8065; // @[Bitwise.scala 50:65:@7460.4]
  wire  _T_8066; // @[Bitwise.scala 50:65:@7461.4]
  wire  _T_8067; // @[Bitwise.scala 50:65:@7462.4]
  wire  _T_8068; // @[Bitwise.scala 50:65:@7463.4]
  wire  _T_8069; // @[Bitwise.scala 50:65:@7464.4]
  wire  _T_8070; // @[Bitwise.scala 50:65:@7465.4]
  wire  _T_8071; // @[Bitwise.scala 50:65:@7466.4]
  wire  _T_8072; // @[Bitwise.scala 50:65:@7467.4]
  wire  _T_8073; // @[Bitwise.scala 50:65:@7468.4]
  wire  _T_8074; // @[Bitwise.scala 50:65:@7469.4]
  wire  _T_8075; // @[Bitwise.scala 50:65:@7470.4]
  wire  _T_8076; // @[Bitwise.scala 50:65:@7471.4]
  wire  _T_8077; // @[Bitwise.scala 50:65:@7472.4]
  wire  _T_8078; // @[Bitwise.scala 50:65:@7473.4]
  wire  _T_8079; // @[Bitwise.scala 50:65:@7474.4]
  wire  _T_8080; // @[Bitwise.scala 50:65:@7475.4]
  wire [1:0] _T_8081; // @[Bitwise.scala 48:55:@7476.4]
  wire [1:0] _GEN_976; // @[Bitwise.scala 48:55:@7477.4]
  wire [2:0] _T_8082; // @[Bitwise.scala 48:55:@7477.4]
  wire [1:0] _T_8083; // @[Bitwise.scala 48:55:@7478.4]
  wire [1:0] _T_8084; // @[Bitwise.scala 48:55:@7479.4]
  wire [2:0] _T_8085; // @[Bitwise.scala 48:55:@7480.4]
  wire [3:0] _T_8086; // @[Bitwise.scala 48:55:@7481.4]
  wire [1:0] _T_8087; // @[Bitwise.scala 48:55:@7482.4]
  wire [1:0] _GEN_977; // @[Bitwise.scala 48:55:@7483.4]
  wire [2:0] _T_8088; // @[Bitwise.scala 48:55:@7483.4]
  wire [1:0] _T_8089; // @[Bitwise.scala 48:55:@7484.4]
  wire [1:0] _T_8090; // @[Bitwise.scala 48:55:@7485.4]
  wire [2:0] _T_8091; // @[Bitwise.scala 48:55:@7486.4]
  wire [3:0] _T_8092; // @[Bitwise.scala 48:55:@7487.4]
  wire [4:0] _T_8093; // @[Bitwise.scala 48:55:@7488.4]
  wire [1:0] _T_8094; // @[Bitwise.scala 48:55:@7489.4]
  wire [1:0] _GEN_978; // @[Bitwise.scala 48:55:@7490.4]
  wire [2:0] _T_8095; // @[Bitwise.scala 48:55:@7490.4]
  wire [1:0] _T_8096; // @[Bitwise.scala 48:55:@7491.4]
  wire [1:0] _T_8097; // @[Bitwise.scala 48:55:@7492.4]
  wire [2:0] _T_8098; // @[Bitwise.scala 48:55:@7493.4]
  wire [3:0] _T_8099; // @[Bitwise.scala 48:55:@7494.4]
  wire [1:0] _T_8100; // @[Bitwise.scala 48:55:@7495.4]
  wire [1:0] _T_8101; // @[Bitwise.scala 48:55:@7496.4]
  wire [2:0] _T_8102; // @[Bitwise.scala 48:55:@7497.4]
  wire [1:0] _T_8103; // @[Bitwise.scala 48:55:@7498.4]
  wire [1:0] _T_8104; // @[Bitwise.scala 48:55:@7499.4]
  wire [2:0] _T_8105; // @[Bitwise.scala 48:55:@7500.4]
  wire [3:0] _T_8106; // @[Bitwise.scala 48:55:@7501.4]
  wire [4:0] _T_8107; // @[Bitwise.scala 48:55:@7502.4]
  wire [5:0] _T_8108; // @[Bitwise.scala 48:55:@7503.4]
  wire [1:0] _T_8109; // @[Bitwise.scala 48:55:@7504.4]
  wire [1:0] _GEN_979; // @[Bitwise.scala 48:55:@7505.4]
  wire [2:0] _T_8110; // @[Bitwise.scala 48:55:@7505.4]
  wire [1:0] _T_8111; // @[Bitwise.scala 48:55:@7506.4]
  wire [1:0] _T_8112; // @[Bitwise.scala 48:55:@7507.4]
  wire [2:0] _T_8113; // @[Bitwise.scala 48:55:@7508.4]
  wire [3:0] _T_8114; // @[Bitwise.scala 48:55:@7509.4]
  wire [1:0] _T_8115; // @[Bitwise.scala 48:55:@7510.4]
  wire [1:0] _GEN_980; // @[Bitwise.scala 48:55:@7511.4]
  wire [2:0] _T_8116; // @[Bitwise.scala 48:55:@7511.4]
  wire [1:0] _T_8117; // @[Bitwise.scala 48:55:@7512.4]
  wire [1:0] _T_8118; // @[Bitwise.scala 48:55:@7513.4]
  wire [2:0] _T_8119; // @[Bitwise.scala 48:55:@7514.4]
  wire [3:0] _T_8120; // @[Bitwise.scala 48:55:@7515.4]
  wire [4:0] _T_8121; // @[Bitwise.scala 48:55:@7516.4]
  wire [1:0] _T_8122; // @[Bitwise.scala 48:55:@7517.4]
  wire [1:0] _GEN_981; // @[Bitwise.scala 48:55:@7518.4]
  wire [2:0] _T_8123; // @[Bitwise.scala 48:55:@7518.4]
  wire [1:0] _T_8124; // @[Bitwise.scala 48:55:@7519.4]
  wire [1:0] _T_8125; // @[Bitwise.scala 48:55:@7520.4]
  wire [2:0] _T_8126; // @[Bitwise.scala 48:55:@7521.4]
  wire [3:0] _T_8127; // @[Bitwise.scala 48:55:@7522.4]
  wire [1:0] _T_8128; // @[Bitwise.scala 48:55:@7523.4]
  wire [1:0] _T_8129; // @[Bitwise.scala 48:55:@7524.4]
  wire [2:0] _T_8130; // @[Bitwise.scala 48:55:@7525.4]
  wire [1:0] _T_8131; // @[Bitwise.scala 48:55:@7526.4]
  wire [1:0] _T_8132; // @[Bitwise.scala 48:55:@7527.4]
  wire [2:0] _T_8133; // @[Bitwise.scala 48:55:@7528.4]
  wire [3:0] _T_8134; // @[Bitwise.scala 48:55:@7529.4]
  wire [4:0] _T_8135; // @[Bitwise.scala 48:55:@7530.4]
  wire [5:0] _T_8136; // @[Bitwise.scala 48:55:@7531.4]
  wire [6:0] _T_8137; // @[Bitwise.scala 48:55:@7532.4]
  wire [58:0] _T_8201; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7597.4]
  wire  _T_8202; // @[Bitwise.scala 50:65:@7598.4]
  wire  _T_8203; // @[Bitwise.scala 50:65:@7599.4]
  wire  _T_8204; // @[Bitwise.scala 50:65:@7600.4]
  wire  _T_8205; // @[Bitwise.scala 50:65:@7601.4]
  wire  _T_8206; // @[Bitwise.scala 50:65:@7602.4]
  wire  _T_8207; // @[Bitwise.scala 50:65:@7603.4]
  wire  _T_8208; // @[Bitwise.scala 50:65:@7604.4]
  wire  _T_8209; // @[Bitwise.scala 50:65:@7605.4]
  wire  _T_8210; // @[Bitwise.scala 50:65:@7606.4]
  wire  _T_8211; // @[Bitwise.scala 50:65:@7607.4]
  wire  _T_8212; // @[Bitwise.scala 50:65:@7608.4]
  wire  _T_8213; // @[Bitwise.scala 50:65:@7609.4]
  wire  _T_8214; // @[Bitwise.scala 50:65:@7610.4]
  wire  _T_8215; // @[Bitwise.scala 50:65:@7611.4]
  wire  _T_8216; // @[Bitwise.scala 50:65:@7612.4]
  wire  _T_8217; // @[Bitwise.scala 50:65:@7613.4]
  wire  _T_8218; // @[Bitwise.scala 50:65:@7614.4]
  wire  _T_8219; // @[Bitwise.scala 50:65:@7615.4]
  wire  _T_8220; // @[Bitwise.scala 50:65:@7616.4]
  wire  _T_8221; // @[Bitwise.scala 50:65:@7617.4]
  wire  _T_8222; // @[Bitwise.scala 50:65:@7618.4]
  wire  _T_8223; // @[Bitwise.scala 50:65:@7619.4]
  wire  _T_8224; // @[Bitwise.scala 50:65:@7620.4]
  wire  _T_8225; // @[Bitwise.scala 50:65:@7621.4]
  wire  _T_8226; // @[Bitwise.scala 50:65:@7622.4]
  wire  _T_8227; // @[Bitwise.scala 50:65:@7623.4]
  wire  _T_8228; // @[Bitwise.scala 50:65:@7624.4]
  wire  _T_8229; // @[Bitwise.scala 50:65:@7625.4]
  wire  _T_8230; // @[Bitwise.scala 50:65:@7626.4]
  wire  _T_8231; // @[Bitwise.scala 50:65:@7627.4]
  wire  _T_8232; // @[Bitwise.scala 50:65:@7628.4]
  wire  _T_8233; // @[Bitwise.scala 50:65:@7629.4]
  wire  _T_8234; // @[Bitwise.scala 50:65:@7630.4]
  wire  _T_8235; // @[Bitwise.scala 50:65:@7631.4]
  wire  _T_8236; // @[Bitwise.scala 50:65:@7632.4]
  wire  _T_8237; // @[Bitwise.scala 50:65:@7633.4]
  wire  _T_8238; // @[Bitwise.scala 50:65:@7634.4]
  wire  _T_8239; // @[Bitwise.scala 50:65:@7635.4]
  wire  _T_8240; // @[Bitwise.scala 50:65:@7636.4]
  wire  _T_8241; // @[Bitwise.scala 50:65:@7637.4]
  wire  _T_8242; // @[Bitwise.scala 50:65:@7638.4]
  wire  _T_8243; // @[Bitwise.scala 50:65:@7639.4]
  wire  _T_8244; // @[Bitwise.scala 50:65:@7640.4]
  wire  _T_8245; // @[Bitwise.scala 50:65:@7641.4]
  wire  _T_8246; // @[Bitwise.scala 50:65:@7642.4]
  wire  _T_8247; // @[Bitwise.scala 50:65:@7643.4]
  wire  _T_8248; // @[Bitwise.scala 50:65:@7644.4]
  wire  _T_8249; // @[Bitwise.scala 50:65:@7645.4]
  wire  _T_8250; // @[Bitwise.scala 50:65:@7646.4]
  wire  _T_8251; // @[Bitwise.scala 50:65:@7647.4]
  wire  _T_8252; // @[Bitwise.scala 50:65:@7648.4]
  wire  _T_8253; // @[Bitwise.scala 50:65:@7649.4]
  wire  _T_8254; // @[Bitwise.scala 50:65:@7650.4]
  wire  _T_8255; // @[Bitwise.scala 50:65:@7651.4]
  wire  _T_8256; // @[Bitwise.scala 50:65:@7652.4]
  wire  _T_8257; // @[Bitwise.scala 50:65:@7653.4]
  wire  _T_8258; // @[Bitwise.scala 50:65:@7654.4]
  wire  _T_8259; // @[Bitwise.scala 50:65:@7655.4]
  wire  _T_8260; // @[Bitwise.scala 50:65:@7656.4]
  wire [1:0] _T_8261; // @[Bitwise.scala 48:55:@7657.4]
  wire [1:0] _GEN_982; // @[Bitwise.scala 48:55:@7658.4]
  wire [2:0] _T_8262; // @[Bitwise.scala 48:55:@7658.4]
  wire [1:0] _T_8263; // @[Bitwise.scala 48:55:@7659.4]
  wire [1:0] _T_8264; // @[Bitwise.scala 48:55:@7660.4]
  wire [2:0] _T_8265; // @[Bitwise.scala 48:55:@7661.4]
  wire [3:0] _T_8266; // @[Bitwise.scala 48:55:@7662.4]
  wire [1:0] _T_8267; // @[Bitwise.scala 48:55:@7663.4]
  wire [1:0] _GEN_983; // @[Bitwise.scala 48:55:@7664.4]
  wire [2:0] _T_8268; // @[Bitwise.scala 48:55:@7664.4]
  wire [1:0] _T_8269; // @[Bitwise.scala 48:55:@7665.4]
  wire [1:0] _T_8270; // @[Bitwise.scala 48:55:@7666.4]
  wire [2:0] _T_8271; // @[Bitwise.scala 48:55:@7667.4]
  wire [3:0] _T_8272; // @[Bitwise.scala 48:55:@7668.4]
  wire [4:0] _T_8273; // @[Bitwise.scala 48:55:@7669.4]
  wire [1:0] _T_8274; // @[Bitwise.scala 48:55:@7670.4]
  wire [1:0] _GEN_984; // @[Bitwise.scala 48:55:@7671.4]
  wire [2:0] _T_8275; // @[Bitwise.scala 48:55:@7671.4]
  wire [1:0] _T_8276; // @[Bitwise.scala 48:55:@7672.4]
  wire [1:0] _T_8277; // @[Bitwise.scala 48:55:@7673.4]
  wire [2:0] _T_8278; // @[Bitwise.scala 48:55:@7674.4]
  wire [3:0] _T_8279; // @[Bitwise.scala 48:55:@7675.4]
  wire [1:0] _T_8280; // @[Bitwise.scala 48:55:@7676.4]
  wire [1:0] _T_8281; // @[Bitwise.scala 48:55:@7677.4]
  wire [2:0] _T_8282; // @[Bitwise.scala 48:55:@7678.4]
  wire [1:0] _T_8283; // @[Bitwise.scala 48:55:@7679.4]
  wire [1:0] _T_8284; // @[Bitwise.scala 48:55:@7680.4]
  wire [2:0] _T_8285; // @[Bitwise.scala 48:55:@7681.4]
  wire [3:0] _T_8286; // @[Bitwise.scala 48:55:@7682.4]
  wire [4:0] _T_8287; // @[Bitwise.scala 48:55:@7683.4]
  wire [5:0] _T_8288; // @[Bitwise.scala 48:55:@7684.4]
  wire [1:0] _T_8289; // @[Bitwise.scala 48:55:@7685.4]
  wire [1:0] _GEN_985; // @[Bitwise.scala 48:55:@7686.4]
  wire [2:0] _T_8290; // @[Bitwise.scala 48:55:@7686.4]
  wire [1:0] _T_8291; // @[Bitwise.scala 48:55:@7687.4]
  wire [1:0] _T_8292; // @[Bitwise.scala 48:55:@7688.4]
  wire [2:0] _T_8293; // @[Bitwise.scala 48:55:@7689.4]
  wire [3:0] _T_8294; // @[Bitwise.scala 48:55:@7690.4]
  wire [1:0] _T_8295; // @[Bitwise.scala 48:55:@7691.4]
  wire [1:0] _T_8296; // @[Bitwise.scala 48:55:@7692.4]
  wire [2:0] _T_8297; // @[Bitwise.scala 48:55:@7693.4]
  wire [1:0] _T_8298; // @[Bitwise.scala 48:55:@7694.4]
  wire [1:0] _T_8299; // @[Bitwise.scala 48:55:@7695.4]
  wire [2:0] _T_8300; // @[Bitwise.scala 48:55:@7696.4]
  wire [3:0] _T_8301; // @[Bitwise.scala 48:55:@7697.4]
  wire [4:0] _T_8302; // @[Bitwise.scala 48:55:@7698.4]
  wire [1:0] _T_8303; // @[Bitwise.scala 48:55:@7699.4]
  wire [1:0] _GEN_986; // @[Bitwise.scala 48:55:@7700.4]
  wire [2:0] _T_8304; // @[Bitwise.scala 48:55:@7700.4]
  wire [1:0] _T_8305; // @[Bitwise.scala 48:55:@7701.4]
  wire [1:0] _T_8306; // @[Bitwise.scala 48:55:@7702.4]
  wire [2:0] _T_8307; // @[Bitwise.scala 48:55:@7703.4]
  wire [3:0] _T_8308; // @[Bitwise.scala 48:55:@7704.4]
  wire [1:0] _T_8309; // @[Bitwise.scala 48:55:@7705.4]
  wire [1:0] _T_8310; // @[Bitwise.scala 48:55:@7706.4]
  wire [2:0] _T_8311; // @[Bitwise.scala 48:55:@7707.4]
  wire [1:0] _T_8312; // @[Bitwise.scala 48:55:@7708.4]
  wire [1:0] _T_8313; // @[Bitwise.scala 48:55:@7709.4]
  wire [2:0] _T_8314; // @[Bitwise.scala 48:55:@7710.4]
  wire [3:0] _T_8315; // @[Bitwise.scala 48:55:@7711.4]
  wire [4:0] _T_8316; // @[Bitwise.scala 48:55:@7712.4]
  wire [5:0] _T_8317; // @[Bitwise.scala 48:55:@7713.4]
  wire [6:0] _T_8318; // @[Bitwise.scala 48:55:@7714.4]
  wire [59:0] _T_8382; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7779.4]
  wire  _T_8383; // @[Bitwise.scala 50:65:@7780.4]
  wire  _T_8384; // @[Bitwise.scala 50:65:@7781.4]
  wire  _T_8385; // @[Bitwise.scala 50:65:@7782.4]
  wire  _T_8386; // @[Bitwise.scala 50:65:@7783.4]
  wire  _T_8387; // @[Bitwise.scala 50:65:@7784.4]
  wire  _T_8388; // @[Bitwise.scala 50:65:@7785.4]
  wire  _T_8389; // @[Bitwise.scala 50:65:@7786.4]
  wire  _T_8390; // @[Bitwise.scala 50:65:@7787.4]
  wire  _T_8391; // @[Bitwise.scala 50:65:@7788.4]
  wire  _T_8392; // @[Bitwise.scala 50:65:@7789.4]
  wire  _T_8393; // @[Bitwise.scala 50:65:@7790.4]
  wire  _T_8394; // @[Bitwise.scala 50:65:@7791.4]
  wire  _T_8395; // @[Bitwise.scala 50:65:@7792.4]
  wire  _T_8396; // @[Bitwise.scala 50:65:@7793.4]
  wire  _T_8397; // @[Bitwise.scala 50:65:@7794.4]
  wire  _T_8398; // @[Bitwise.scala 50:65:@7795.4]
  wire  _T_8399; // @[Bitwise.scala 50:65:@7796.4]
  wire  _T_8400; // @[Bitwise.scala 50:65:@7797.4]
  wire  _T_8401; // @[Bitwise.scala 50:65:@7798.4]
  wire  _T_8402; // @[Bitwise.scala 50:65:@7799.4]
  wire  _T_8403; // @[Bitwise.scala 50:65:@7800.4]
  wire  _T_8404; // @[Bitwise.scala 50:65:@7801.4]
  wire  _T_8405; // @[Bitwise.scala 50:65:@7802.4]
  wire  _T_8406; // @[Bitwise.scala 50:65:@7803.4]
  wire  _T_8407; // @[Bitwise.scala 50:65:@7804.4]
  wire  _T_8408; // @[Bitwise.scala 50:65:@7805.4]
  wire  _T_8409; // @[Bitwise.scala 50:65:@7806.4]
  wire  _T_8410; // @[Bitwise.scala 50:65:@7807.4]
  wire  _T_8411; // @[Bitwise.scala 50:65:@7808.4]
  wire  _T_8412; // @[Bitwise.scala 50:65:@7809.4]
  wire  _T_8413; // @[Bitwise.scala 50:65:@7810.4]
  wire  _T_8414; // @[Bitwise.scala 50:65:@7811.4]
  wire  _T_8415; // @[Bitwise.scala 50:65:@7812.4]
  wire  _T_8416; // @[Bitwise.scala 50:65:@7813.4]
  wire  _T_8417; // @[Bitwise.scala 50:65:@7814.4]
  wire  _T_8418; // @[Bitwise.scala 50:65:@7815.4]
  wire  _T_8419; // @[Bitwise.scala 50:65:@7816.4]
  wire  _T_8420; // @[Bitwise.scala 50:65:@7817.4]
  wire  _T_8421; // @[Bitwise.scala 50:65:@7818.4]
  wire  _T_8422; // @[Bitwise.scala 50:65:@7819.4]
  wire  _T_8423; // @[Bitwise.scala 50:65:@7820.4]
  wire  _T_8424; // @[Bitwise.scala 50:65:@7821.4]
  wire  _T_8425; // @[Bitwise.scala 50:65:@7822.4]
  wire  _T_8426; // @[Bitwise.scala 50:65:@7823.4]
  wire  _T_8427; // @[Bitwise.scala 50:65:@7824.4]
  wire  _T_8428; // @[Bitwise.scala 50:65:@7825.4]
  wire  _T_8429; // @[Bitwise.scala 50:65:@7826.4]
  wire  _T_8430; // @[Bitwise.scala 50:65:@7827.4]
  wire  _T_8431; // @[Bitwise.scala 50:65:@7828.4]
  wire  _T_8432; // @[Bitwise.scala 50:65:@7829.4]
  wire  _T_8433; // @[Bitwise.scala 50:65:@7830.4]
  wire  _T_8434; // @[Bitwise.scala 50:65:@7831.4]
  wire  _T_8435; // @[Bitwise.scala 50:65:@7832.4]
  wire  _T_8436; // @[Bitwise.scala 50:65:@7833.4]
  wire  _T_8437; // @[Bitwise.scala 50:65:@7834.4]
  wire  _T_8438; // @[Bitwise.scala 50:65:@7835.4]
  wire  _T_8439; // @[Bitwise.scala 50:65:@7836.4]
  wire  _T_8440; // @[Bitwise.scala 50:65:@7837.4]
  wire  _T_8441; // @[Bitwise.scala 50:65:@7838.4]
  wire  _T_8442; // @[Bitwise.scala 50:65:@7839.4]
  wire [1:0] _T_8443; // @[Bitwise.scala 48:55:@7840.4]
  wire [1:0] _GEN_987; // @[Bitwise.scala 48:55:@7841.4]
  wire [2:0] _T_8444; // @[Bitwise.scala 48:55:@7841.4]
  wire [1:0] _T_8445; // @[Bitwise.scala 48:55:@7842.4]
  wire [1:0] _T_8446; // @[Bitwise.scala 48:55:@7843.4]
  wire [2:0] _T_8447; // @[Bitwise.scala 48:55:@7844.4]
  wire [3:0] _T_8448; // @[Bitwise.scala 48:55:@7845.4]
  wire [1:0] _T_8449; // @[Bitwise.scala 48:55:@7846.4]
  wire [1:0] _T_8450; // @[Bitwise.scala 48:55:@7847.4]
  wire [2:0] _T_8451; // @[Bitwise.scala 48:55:@7848.4]
  wire [1:0] _T_8452; // @[Bitwise.scala 48:55:@7849.4]
  wire [1:0] _T_8453; // @[Bitwise.scala 48:55:@7850.4]
  wire [2:0] _T_8454; // @[Bitwise.scala 48:55:@7851.4]
  wire [3:0] _T_8455; // @[Bitwise.scala 48:55:@7852.4]
  wire [4:0] _T_8456; // @[Bitwise.scala 48:55:@7853.4]
  wire [1:0] _T_8457; // @[Bitwise.scala 48:55:@7854.4]
  wire [1:0] _GEN_988; // @[Bitwise.scala 48:55:@7855.4]
  wire [2:0] _T_8458; // @[Bitwise.scala 48:55:@7855.4]
  wire [1:0] _T_8459; // @[Bitwise.scala 48:55:@7856.4]
  wire [1:0] _T_8460; // @[Bitwise.scala 48:55:@7857.4]
  wire [2:0] _T_8461; // @[Bitwise.scala 48:55:@7858.4]
  wire [3:0] _T_8462; // @[Bitwise.scala 48:55:@7859.4]
  wire [1:0] _T_8463; // @[Bitwise.scala 48:55:@7860.4]
  wire [1:0] _T_8464; // @[Bitwise.scala 48:55:@7861.4]
  wire [2:0] _T_8465; // @[Bitwise.scala 48:55:@7862.4]
  wire [1:0] _T_8466; // @[Bitwise.scala 48:55:@7863.4]
  wire [1:0] _T_8467; // @[Bitwise.scala 48:55:@7864.4]
  wire [2:0] _T_8468; // @[Bitwise.scala 48:55:@7865.4]
  wire [3:0] _T_8469; // @[Bitwise.scala 48:55:@7866.4]
  wire [4:0] _T_8470; // @[Bitwise.scala 48:55:@7867.4]
  wire [5:0] _T_8471; // @[Bitwise.scala 48:55:@7868.4]
  wire [1:0] _T_8472; // @[Bitwise.scala 48:55:@7869.4]
  wire [1:0] _GEN_989; // @[Bitwise.scala 48:55:@7870.4]
  wire [2:0] _T_8473; // @[Bitwise.scala 48:55:@7870.4]
  wire [1:0] _T_8474; // @[Bitwise.scala 48:55:@7871.4]
  wire [1:0] _T_8475; // @[Bitwise.scala 48:55:@7872.4]
  wire [2:0] _T_8476; // @[Bitwise.scala 48:55:@7873.4]
  wire [3:0] _T_8477; // @[Bitwise.scala 48:55:@7874.4]
  wire [1:0] _T_8478; // @[Bitwise.scala 48:55:@7875.4]
  wire [1:0] _T_8479; // @[Bitwise.scala 48:55:@7876.4]
  wire [2:0] _T_8480; // @[Bitwise.scala 48:55:@7877.4]
  wire [1:0] _T_8481; // @[Bitwise.scala 48:55:@7878.4]
  wire [1:0] _T_8482; // @[Bitwise.scala 48:55:@7879.4]
  wire [2:0] _T_8483; // @[Bitwise.scala 48:55:@7880.4]
  wire [3:0] _T_8484; // @[Bitwise.scala 48:55:@7881.4]
  wire [4:0] _T_8485; // @[Bitwise.scala 48:55:@7882.4]
  wire [1:0] _T_8486; // @[Bitwise.scala 48:55:@7883.4]
  wire [1:0] _GEN_990; // @[Bitwise.scala 48:55:@7884.4]
  wire [2:0] _T_8487; // @[Bitwise.scala 48:55:@7884.4]
  wire [1:0] _T_8488; // @[Bitwise.scala 48:55:@7885.4]
  wire [1:0] _T_8489; // @[Bitwise.scala 48:55:@7886.4]
  wire [2:0] _T_8490; // @[Bitwise.scala 48:55:@7887.4]
  wire [3:0] _T_8491; // @[Bitwise.scala 48:55:@7888.4]
  wire [1:0] _T_8492; // @[Bitwise.scala 48:55:@7889.4]
  wire [1:0] _T_8493; // @[Bitwise.scala 48:55:@7890.4]
  wire [2:0] _T_8494; // @[Bitwise.scala 48:55:@7891.4]
  wire [1:0] _T_8495; // @[Bitwise.scala 48:55:@7892.4]
  wire [1:0] _T_8496; // @[Bitwise.scala 48:55:@7893.4]
  wire [2:0] _T_8497; // @[Bitwise.scala 48:55:@7894.4]
  wire [3:0] _T_8498; // @[Bitwise.scala 48:55:@7895.4]
  wire [4:0] _T_8499; // @[Bitwise.scala 48:55:@7896.4]
  wire [5:0] _T_8500; // @[Bitwise.scala 48:55:@7897.4]
  wire [6:0] _T_8501; // @[Bitwise.scala 48:55:@7898.4]
  wire [60:0] _T_8565; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7963.4]
  wire  _T_8566; // @[Bitwise.scala 50:65:@7964.4]
  wire  _T_8567; // @[Bitwise.scala 50:65:@7965.4]
  wire  _T_8568; // @[Bitwise.scala 50:65:@7966.4]
  wire  _T_8569; // @[Bitwise.scala 50:65:@7967.4]
  wire  _T_8570; // @[Bitwise.scala 50:65:@7968.4]
  wire  _T_8571; // @[Bitwise.scala 50:65:@7969.4]
  wire  _T_8572; // @[Bitwise.scala 50:65:@7970.4]
  wire  _T_8573; // @[Bitwise.scala 50:65:@7971.4]
  wire  _T_8574; // @[Bitwise.scala 50:65:@7972.4]
  wire  _T_8575; // @[Bitwise.scala 50:65:@7973.4]
  wire  _T_8576; // @[Bitwise.scala 50:65:@7974.4]
  wire  _T_8577; // @[Bitwise.scala 50:65:@7975.4]
  wire  _T_8578; // @[Bitwise.scala 50:65:@7976.4]
  wire  _T_8579; // @[Bitwise.scala 50:65:@7977.4]
  wire  _T_8580; // @[Bitwise.scala 50:65:@7978.4]
  wire  _T_8581; // @[Bitwise.scala 50:65:@7979.4]
  wire  _T_8582; // @[Bitwise.scala 50:65:@7980.4]
  wire  _T_8583; // @[Bitwise.scala 50:65:@7981.4]
  wire  _T_8584; // @[Bitwise.scala 50:65:@7982.4]
  wire  _T_8585; // @[Bitwise.scala 50:65:@7983.4]
  wire  _T_8586; // @[Bitwise.scala 50:65:@7984.4]
  wire  _T_8587; // @[Bitwise.scala 50:65:@7985.4]
  wire  _T_8588; // @[Bitwise.scala 50:65:@7986.4]
  wire  _T_8589; // @[Bitwise.scala 50:65:@7987.4]
  wire  _T_8590; // @[Bitwise.scala 50:65:@7988.4]
  wire  _T_8591; // @[Bitwise.scala 50:65:@7989.4]
  wire  _T_8592; // @[Bitwise.scala 50:65:@7990.4]
  wire  _T_8593; // @[Bitwise.scala 50:65:@7991.4]
  wire  _T_8594; // @[Bitwise.scala 50:65:@7992.4]
  wire  _T_8595; // @[Bitwise.scala 50:65:@7993.4]
  wire  _T_8596; // @[Bitwise.scala 50:65:@7994.4]
  wire  _T_8597; // @[Bitwise.scala 50:65:@7995.4]
  wire  _T_8598; // @[Bitwise.scala 50:65:@7996.4]
  wire  _T_8599; // @[Bitwise.scala 50:65:@7997.4]
  wire  _T_8600; // @[Bitwise.scala 50:65:@7998.4]
  wire  _T_8601; // @[Bitwise.scala 50:65:@7999.4]
  wire  _T_8602; // @[Bitwise.scala 50:65:@8000.4]
  wire  _T_8603; // @[Bitwise.scala 50:65:@8001.4]
  wire  _T_8604; // @[Bitwise.scala 50:65:@8002.4]
  wire  _T_8605; // @[Bitwise.scala 50:65:@8003.4]
  wire  _T_8606; // @[Bitwise.scala 50:65:@8004.4]
  wire  _T_8607; // @[Bitwise.scala 50:65:@8005.4]
  wire  _T_8608; // @[Bitwise.scala 50:65:@8006.4]
  wire  _T_8609; // @[Bitwise.scala 50:65:@8007.4]
  wire  _T_8610; // @[Bitwise.scala 50:65:@8008.4]
  wire  _T_8611; // @[Bitwise.scala 50:65:@8009.4]
  wire  _T_8612; // @[Bitwise.scala 50:65:@8010.4]
  wire  _T_8613; // @[Bitwise.scala 50:65:@8011.4]
  wire  _T_8614; // @[Bitwise.scala 50:65:@8012.4]
  wire  _T_8615; // @[Bitwise.scala 50:65:@8013.4]
  wire  _T_8616; // @[Bitwise.scala 50:65:@8014.4]
  wire  _T_8617; // @[Bitwise.scala 50:65:@8015.4]
  wire  _T_8618; // @[Bitwise.scala 50:65:@8016.4]
  wire  _T_8619; // @[Bitwise.scala 50:65:@8017.4]
  wire  _T_8620; // @[Bitwise.scala 50:65:@8018.4]
  wire  _T_8621; // @[Bitwise.scala 50:65:@8019.4]
  wire  _T_8622; // @[Bitwise.scala 50:65:@8020.4]
  wire  _T_8623; // @[Bitwise.scala 50:65:@8021.4]
  wire  _T_8624; // @[Bitwise.scala 50:65:@8022.4]
  wire  _T_8625; // @[Bitwise.scala 50:65:@8023.4]
  wire  _T_8626; // @[Bitwise.scala 50:65:@8024.4]
  wire [1:0] _T_8627; // @[Bitwise.scala 48:55:@8025.4]
  wire [1:0] _GEN_991; // @[Bitwise.scala 48:55:@8026.4]
  wire [2:0] _T_8628; // @[Bitwise.scala 48:55:@8026.4]
  wire [1:0] _T_8629; // @[Bitwise.scala 48:55:@8027.4]
  wire [1:0] _T_8630; // @[Bitwise.scala 48:55:@8028.4]
  wire [2:0] _T_8631; // @[Bitwise.scala 48:55:@8029.4]
  wire [3:0] _T_8632; // @[Bitwise.scala 48:55:@8030.4]
  wire [1:0] _T_8633; // @[Bitwise.scala 48:55:@8031.4]
  wire [1:0] _T_8634; // @[Bitwise.scala 48:55:@8032.4]
  wire [2:0] _T_8635; // @[Bitwise.scala 48:55:@8033.4]
  wire [1:0] _T_8636; // @[Bitwise.scala 48:55:@8034.4]
  wire [1:0] _T_8637; // @[Bitwise.scala 48:55:@8035.4]
  wire [2:0] _T_8638; // @[Bitwise.scala 48:55:@8036.4]
  wire [3:0] _T_8639; // @[Bitwise.scala 48:55:@8037.4]
  wire [4:0] _T_8640; // @[Bitwise.scala 48:55:@8038.4]
  wire [1:0] _T_8641; // @[Bitwise.scala 48:55:@8039.4]
  wire [1:0] _GEN_992; // @[Bitwise.scala 48:55:@8040.4]
  wire [2:0] _T_8642; // @[Bitwise.scala 48:55:@8040.4]
  wire [1:0] _T_8643; // @[Bitwise.scala 48:55:@8041.4]
  wire [1:0] _T_8644; // @[Bitwise.scala 48:55:@8042.4]
  wire [2:0] _T_8645; // @[Bitwise.scala 48:55:@8043.4]
  wire [3:0] _T_8646; // @[Bitwise.scala 48:55:@8044.4]
  wire [1:0] _T_8647; // @[Bitwise.scala 48:55:@8045.4]
  wire [1:0] _T_8648; // @[Bitwise.scala 48:55:@8046.4]
  wire [2:0] _T_8649; // @[Bitwise.scala 48:55:@8047.4]
  wire [1:0] _T_8650; // @[Bitwise.scala 48:55:@8048.4]
  wire [1:0] _T_8651; // @[Bitwise.scala 48:55:@8049.4]
  wire [2:0] _T_8652; // @[Bitwise.scala 48:55:@8050.4]
  wire [3:0] _T_8653; // @[Bitwise.scala 48:55:@8051.4]
  wire [4:0] _T_8654; // @[Bitwise.scala 48:55:@8052.4]
  wire [5:0] _T_8655; // @[Bitwise.scala 48:55:@8053.4]
  wire [1:0] _T_8656; // @[Bitwise.scala 48:55:@8054.4]
  wire [1:0] _GEN_993; // @[Bitwise.scala 48:55:@8055.4]
  wire [2:0] _T_8657; // @[Bitwise.scala 48:55:@8055.4]
  wire [1:0] _T_8658; // @[Bitwise.scala 48:55:@8056.4]
  wire [1:0] _T_8659; // @[Bitwise.scala 48:55:@8057.4]
  wire [2:0] _T_8660; // @[Bitwise.scala 48:55:@8058.4]
  wire [3:0] _T_8661; // @[Bitwise.scala 48:55:@8059.4]
  wire [1:0] _T_8662; // @[Bitwise.scala 48:55:@8060.4]
  wire [1:0] _T_8663; // @[Bitwise.scala 48:55:@8061.4]
  wire [2:0] _T_8664; // @[Bitwise.scala 48:55:@8062.4]
  wire [1:0] _T_8665; // @[Bitwise.scala 48:55:@8063.4]
  wire [1:0] _T_8666; // @[Bitwise.scala 48:55:@8064.4]
  wire [2:0] _T_8667; // @[Bitwise.scala 48:55:@8065.4]
  wire [3:0] _T_8668; // @[Bitwise.scala 48:55:@8066.4]
  wire [4:0] _T_8669; // @[Bitwise.scala 48:55:@8067.4]
  wire [1:0] _T_8670; // @[Bitwise.scala 48:55:@8068.4]
  wire [1:0] _T_8671; // @[Bitwise.scala 48:55:@8069.4]
  wire [2:0] _T_8672; // @[Bitwise.scala 48:55:@8070.4]
  wire [1:0] _T_8673; // @[Bitwise.scala 48:55:@8071.4]
  wire [1:0] _T_8674; // @[Bitwise.scala 48:55:@8072.4]
  wire [2:0] _T_8675; // @[Bitwise.scala 48:55:@8073.4]
  wire [3:0] _T_8676; // @[Bitwise.scala 48:55:@8074.4]
  wire [1:0] _T_8677; // @[Bitwise.scala 48:55:@8075.4]
  wire [1:0] _T_8678; // @[Bitwise.scala 48:55:@8076.4]
  wire [2:0] _T_8679; // @[Bitwise.scala 48:55:@8077.4]
  wire [1:0] _T_8680; // @[Bitwise.scala 48:55:@8078.4]
  wire [1:0] _T_8681; // @[Bitwise.scala 48:55:@8079.4]
  wire [2:0] _T_8682; // @[Bitwise.scala 48:55:@8080.4]
  wire [3:0] _T_8683; // @[Bitwise.scala 48:55:@8081.4]
  wire [4:0] _T_8684; // @[Bitwise.scala 48:55:@8082.4]
  wire [5:0] _T_8685; // @[Bitwise.scala 48:55:@8083.4]
  wire [6:0] _T_8686; // @[Bitwise.scala 48:55:@8084.4]
  wire [61:0] _T_8750; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@8149.4]
  wire  _T_8751; // @[Bitwise.scala 50:65:@8150.4]
  wire  _T_8752; // @[Bitwise.scala 50:65:@8151.4]
  wire  _T_8753; // @[Bitwise.scala 50:65:@8152.4]
  wire  _T_8754; // @[Bitwise.scala 50:65:@8153.4]
  wire  _T_8755; // @[Bitwise.scala 50:65:@8154.4]
  wire  _T_8756; // @[Bitwise.scala 50:65:@8155.4]
  wire  _T_8757; // @[Bitwise.scala 50:65:@8156.4]
  wire  _T_8758; // @[Bitwise.scala 50:65:@8157.4]
  wire  _T_8759; // @[Bitwise.scala 50:65:@8158.4]
  wire  _T_8760; // @[Bitwise.scala 50:65:@8159.4]
  wire  _T_8761; // @[Bitwise.scala 50:65:@8160.4]
  wire  _T_8762; // @[Bitwise.scala 50:65:@8161.4]
  wire  _T_8763; // @[Bitwise.scala 50:65:@8162.4]
  wire  _T_8764; // @[Bitwise.scala 50:65:@8163.4]
  wire  _T_8765; // @[Bitwise.scala 50:65:@8164.4]
  wire  _T_8766; // @[Bitwise.scala 50:65:@8165.4]
  wire  _T_8767; // @[Bitwise.scala 50:65:@8166.4]
  wire  _T_8768; // @[Bitwise.scala 50:65:@8167.4]
  wire  _T_8769; // @[Bitwise.scala 50:65:@8168.4]
  wire  _T_8770; // @[Bitwise.scala 50:65:@8169.4]
  wire  _T_8771; // @[Bitwise.scala 50:65:@8170.4]
  wire  _T_8772; // @[Bitwise.scala 50:65:@8171.4]
  wire  _T_8773; // @[Bitwise.scala 50:65:@8172.4]
  wire  _T_8774; // @[Bitwise.scala 50:65:@8173.4]
  wire  _T_8775; // @[Bitwise.scala 50:65:@8174.4]
  wire  _T_8776; // @[Bitwise.scala 50:65:@8175.4]
  wire  _T_8777; // @[Bitwise.scala 50:65:@8176.4]
  wire  _T_8778; // @[Bitwise.scala 50:65:@8177.4]
  wire  _T_8779; // @[Bitwise.scala 50:65:@8178.4]
  wire  _T_8780; // @[Bitwise.scala 50:65:@8179.4]
  wire  _T_8781; // @[Bitwise.scala 50:65:@8180.4]
  wire  _T_8782; // @[Bitwise.scala 50:65:@8181.4]
  wire  _T_8783; // @[Bitwise.scala 50:65:@8182.4]
  wire  _T_8784; // @[Bitwise.scala 50:65:@8183.4]
  wire  _T_8785; // @[Bitwise.scala 50:65:@8184.4]
  wire  _T_8786; // @[Bitwise.scala 50:65:@8185.4]
  wire  _T_8787; // @[Bitwise.scala 50:65:@8186.4]
  wire  _T_8788; // @[Bitwise.scala 50:65:@8187.4]
  wire  _T_8789; // @[Bitwise.scala 50:65:@8188.4]
  wire  _T_8790; // @[Bitwise.scala 50:65:@8189.4]
  wire  _T_8791; // @[Bitwise.scala 50:65:@8190.4]
  wire  _T_8792; // @[Bitwise.scala 50:65:@8191.4]
  wire  _T_8793; // @[Bitwise.scala 50:65:@8192.4]
  wire  _T_8794; // @[Bitwise.scala 50:65:@8193.4]
  wire  _T_8795; // @[Bitwise.scala 50:65:@8194.4]
  wire  _T_8796; // @[Bitwise.scala 50:65:@8195.4]
  wire  _T_8797; // @[Bitwise.scala 50:65:@8196.4]
  wire  _T_8798; // @[Bitwise.scala 50:65:@8197.4]
  wire  _T_8799; // @[Bitwise.scala 50:65:@8198.4]
  wire  _T_8800; // @[Bitwise.scala 50:65:@8199.4]
  wire  _T_8801; // @[Bitwise.scala 50:65:@8200.4]
  wire  _T_8802; // @[Bitwise.scala 50:65:@8201.4]
  wire  _T_8803; // @[Bitwise.scala 50:65:@8202.4]
  wire  _T_8804; // @[Bitwise.scala 50:65:@8203.4]
  wire  _T_8805; // @[Bitwise.scala 50:65:@8204.4]
  wire  _T_8806; // @[Bitwise.scala 50:65:@8205.4]
  wire  _T_8807; // @[Bitwise.scala 50:65:@8206.4]
  wire  _T_8808; // @[Bitwise.scala 50:65:@8207.4]
  wire  _T_8809; // @[Bitwise.scala 50:65:@8208.4]
  wire  _T_8810; // @[Bitwise.scala 50:65:@8209.4]
  wire  _T_8811; // @[Bitwise.scala 50:65:@8210.4]
  wire  _T_8812; // @[Bitwise.scala 50:65:@8211.4]
  wire [1:0] _T_8813; // @[Bitwise.scala 48:55:@8212.4]
  wire [1:0] _GEN_994; // @[Bitwise.scala 48:55:@8213.4]
  wire [2:0] _T_8814; // @[Bitwise.scala 48:55:@8213.4]
  wire [1:0] _T_8815; // @[Bitwise.scala 48:55:@8214.4]
  wire [1:0] _T_8816; // @[Bitwise.scala 48:55:@8215.4]
  wire [2:0] _T_8817; // @[Bitwise.scala 48:55:@8216.4]
  wire [3:0] _T_8818; // @[Bitwise.scala 48:55:@8217.4]
  wire [1:0] _T_8819; // @[Bitwise.scala 48:55:@8218.4]
  wire [1:0] _T_8820; // @[Bitwise.scala 48:55:@8219.4]
  wire [2:0] _T_8821; // @[Bitwise.scala 48:55:@8220.4]
  wire [1:0] _T_8822; // @[Bitwise.scala 48:55:@8221.4]
  wire [1:0] _T_8823; // @[Bitwise.scala 48:55:@8222.4]
  wire [2:0] _T_8824; // @[Bitwise.scala 48:55:@8223.4]
  wire [3:0] _T_8825; // @[Bitwise.scala 48:55:@8224.4]
  wire [4:0] _T_8826; // @[Bitwise.scala 48:55:@8225.4]
  wire [1:0] _T_8827; // @[Bitwise.scala 48:55:@8226.4]
  wire [1:0] _T_8828; // @[Bitwise.scala 48:55:@8227.4]
  wire [2:0] _T_8829; // @[Bitwise.scala 48:55:@8228.4]
  wire [1:0] _T_8830; // @[Bitwise.scala 48:55:@8229.4]
  wire [1:0] _T_8831; // @[Bitwise.scala 48:55:@8230.4]
  wire [2:0] _T_8832; // @[Bitwise.scala 48:55:@8231.4]
  wire [3:0] _T_8833; // @[Bitwise.scala 48:55:@8232.4]
  wire [1:0] _T_8834; // @[Bitwise.scala 48:55:@8233.4]
  wire [1:0] _T_8835; // @[Bitwise.scala 48:55:@8234.4]
  wire [2:0] _T_8836; // @[Bitwise.scala 48:55:@8235.4]
  wire [1:0] _T_8837; // @[Bitwise.scala 48:55:@8236.4]
  wire [1:0] _T_8838; // @[Bitwise.scala 48:55:@8237.4]
  wire [2:0] _T_8839; // @[Bitwise.scala 48:55:@8238.4]
  wire [3:0] _T_8840; // @[Bitwise.scala 48:55:@8239.4]
  wire [4:0] _T_8841; // @[Bitwise.scala 48:55:@8240.4]
  wire [5:0] _T_8842; // @[Bitwise.scala 48:55:@8241.4]
  wire [1:0] _T_8843; // @[Bitwise.scala 48:55:@8242.4]
  wire [1:0] _GEN_995; // @[Bitwise.scala 48:55:@8243.4]
  wire [2:0] _T_8844; // @[Bitwise.scala 48:55:@8243.4]
  wire [1:0] _T_8845; // @[Bitwise.scala 48:55:@8244.4]
  wire [1:0] _T_8846; // @[Bitwise.scala 48:55:@8245.4]
  wire [2:0] _T_8847; // @[Bitwise.scala 48:55:@8246.4]
  wire [3:0] _T_8848; // @[Bitwise.scala 48:55:@8247.4]
  wire [1:0] _T_8849; // @[Bitwise.scala 48:55:@8248.4]
  wire [1:0] _T_8850; // @[Bitwise.scala 48:55:@8249.4]
  wire [2:0] _T_8851; // @[Bitwise.scala 48:55:@8250.4]
  wire [1:0] _T_8852; // @[Bitwise.scala 48:55:@8251.4]
  wire [1:0] _T_8853; // @[Bitwise.scala 48:55:@8252.4]
  wire [2:0] _T_8854; // @[Bitwise.scala 48:55:@8253.4]
  wire [3:0] _T_8855; // @[Bitwise.scala 48:55:@8254.4]
  wire [4:0] _T_8856; // @[Bitwise.scala 48:55:@8255.4]
  wire [1:0] _T_8857; // @[Bitwise.scala 48:55:@8256.4]
  wire [1:0] _T_8858; // @[Bitwise.scala 48:55:@8257.4]
  wire [2:0] _T_8859; // @[Bitwise.scala 48:55:@8258.4]
  wire [1:0] _T_8860; // @[Bitwise.scala 48:55:@8259.4]
  wire [1:0] _T_8861; // @[Bitwise.scala 48:55:@8260.4]
  wire [2:0] _T_8862; // @[Bitwise.scala 48:55:@8261.4]
  wire [3:0] _T_8863; // @[Bitwise.scala 48:55:@8262.4]
  wire [1:0] _T_8864; // @[Bitwise.scala 48:55:@8263.4]
  wire [1:0] _T_8865; // @[Bitwise.scala 48:55:@8264.4]
  wire [2:0] _T_8866; // @[Bitwise.scala 48:55:@8265.4]
  wire [1:0] _T_8867; // @[Bitwise.scala 48:55:@8266.4]
  wire [1:0] _T_8868; // @[Bitwise.scala 48:55:@8267.4]
  wire [2:0] _T_8869; // @[Bitwise.scala 48:55:@8268.4]
  wire [3:0] _T_8870; // @[Bitwise.scala 48:55:@8269.4]
  wire [4:0] _T_8871; // @[Bitwise.scala 48:55:@8270.4]
  wire [5:0] _T_8872; // @[Bitwise.scala 48:55:@8271.4]
  wire [6:0] _T_8873; // @[Bitwise.scala 48:55:@8272.4]
  wire [62:0] _T_8937; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@8337.4]
  wire  _T_8938; // @[Bitwise.scala 50:65:@8338.4]
  wire  _T_8939; // @[Bitwise.scala 50:65:@8339.4]
  wire  _T_8940; // @[Bitwise.scala 50:65:@8340.4]
  wire  _T_8941; // @[Bitwise.scala 50:65:@8341.4]
  wire  _T_8942; // @[Bitwise.scala 50:65:@8342.4]
  wire  _T_8943; // @[Bitwise.scala 50:65:@8343.4]
  wire  _T_8944; // @[Bitwise.scala 50:65:@8344.4]
  wire  _T_8945; // @[Bitwise.scala 50:65:@8345.4]
  wire  _T_8946; // @[Bitwise.scala 50:65:@8346.4]
  wire  _T_8947; // @[Bitwise.scala 50:65:@8347.4]
  wire  _T_8948; // @[Bitwise.scala 50:65:@8348.4]
  wire  _T_8949; // @[Bitwise.scala 50:65:@8349.4]
  wire  _T_8950; // @[Bitwise.scala 50:65:@8350.4]
  wire  _T_8951; // @[Bitwise.scala 50:65:@8351.4]
  wire  _T_8952; // @[Bitwise.scala 50:65:@8352.4]
  wire  _T_8953; // @[Bitwise.scala 50:65:@8353.4]
  wire  _T_8954; // @[Bitwise.scala 50:65:@8354.4]
  wire  _T_8955; // @[Bitwise.scala 50:65:@8355.4]
  wire  _T_8956; // @[Bitwise.scala 50:65:@8356.4]
  wire  _T_8957; // @[Bitwise.scala 50:65:@8357.4]
  wire  _T_8958; // @[Bitwise.scala 50:65:@8358.4]
  wire  _T_8959; // @[Bitwise.scala 50:65:@8359.4]
  wire  _T_8960; // @[Bitwise.scala 50:65:@8360.4]
  wire  _T_8961; // @[Bitwise.scala 50:65:@8361.4]
  wire  _T_8962; // @[Bitwise.scala 50:65:@8362.4]
  wire  _T_8963; // @[Bitwise.scala 50:65:@8363.4]
  wire  _T_8964; // @[Bitwise.scala 50:65:@8364.4]
  wire  _T_8965; // @[Bitwise.scala 50:65:@8365.4]
  wire  _T_8966; // @[Bitwise.scala 50:65:@8366.4]
  wire  _T_8967; // @[Bitwise.scala 50:65:@8367.4]
  wire  _T_8968; // @[Bitwise.scala 50:65:@8368.4]
  wire  _T_8969; // @[Bitwise.scala 50:65:@8369.4]
  wire  _T_8970; // @[Bitwise.scala 50:65:@8370.4]
  wire  _T_8971; // @[Bitwise.scala 50:65:@8371.4]
  wire  _T_8972; // @[Bitwise.scala 50:65:@8372.4]
  wire  _T_8973; // @[Bitwise.scala 50:65:@8373.4]
  wire  _T_8974; // @[Bitwise.scala 50:65:@8374.4]
  wire  _T_8975; // @[Bitwise.scala 50:65:@8375.4]
  wire  _T_8976; // @[Bitwise.scala 50:65:@8376.4]
  wire  _T_8977; // @[Bitwise.scala 50:65:@8377.4]
  wire  _T_8978; // @[Bitwise.scala 50:65:@8378.4]
  wire  _T_8979; // @[Bitwise.scala 50:65:@8379.4]
  wire  _T_8980; // @[Bitwise.scala 50:65:@8380.4]
  wire  _T_8981; // @[Bitwise.scala 50:65:@8381.4]
  wire  _T_8982; // @[Bitwise.scala 50:65:@8382.4]
  wire  _T_8983; // @[Bitwise.scala 50:65:@8383.4]
  wire  _T_8984; // @[Bitwise.scala 50:65:@8384.4]
  wire  _T_8985; // @[Bitwise.scala 50:65:@8385.4]
  wire  _T_8986; // @[Bitwise.scala 50:65:@8386.4]
  wire  _T_8987; // @[Bitwise.scala 50:65:@8387.4]
  wire  _T_8988; // @[Bitwise.scala 50:65:@8388.4]
  wire  _T_8989; // @[Bitwise.scala 50:65:@8389.4]
  wire  _T_8990; // @[Bitwise.scala 50:65:@8390.4]
  wire  _T_8991; // @[Bitwise.scala 50:65:@8391.4]
  wire  _T_8992; // @[Bitwise.scala 50:65:@8392.4]
  wire  _T_8993; // @[Bitwise.scala 50:65:@8393.4]
  wire  _T_8994; // @[Bitwise.scala 50:65:@8394.4]
  wire  _T_8995; // @[Bitwise.scala 50:65:@8395.4]
  wire  _T_8996; // @[Bitwise.scala 50:65:@8396.4]
  wire  _T_8997; // @[Bitwise.scala 50:65:@8397.4]
  wire  _T_8998; // @[Bitwise.scala 50:65:@8398.4]
  wire  _T_8999; // @[Bitwise.scala 50:65:@8399.4]
  wire  _T_9000; // @[Bitwise.scala 50:65:@8400.4]
  wire [1:0] _T_9001; // @[Bitwise.scala 48:55:@8401.4]
  wire [1:0] _GEN_996; // @[Bitwise.scala 48:55:@8402.4]
  wire [2:0] _T_9002; // @[Bitwise.scala 48:55:@8402.4]
  wire [1:0] _T_9003; // @[Bitwise.scala 48:55:@8403.4]
  wire [1:0] _T_9004; // @[Bitwise.scala 48:55:@8404.4]
  wire [2:0] _T_9005; // @[Bitwise.scala 48:55:@8405.4]
  wire [3:0] _T_9006; // @[Bitwise.scala 48:55:@8406.4]
  wire [1:0] _T_9007; // @[Bitwise.scala 48:55:@8407.4]
  wire [1:0] _T_9008; // @[Bitwise.scala 48:55:@8408.4]
  wire [2:0] _T_9009; // @[Bitwise.scala 48:55:@8409.4]
  wire [1:0] _T_9010; // @[Bitwise.scala 48:55:@8410.4]
  wire [1:0] _T_9011; // @[Bitwise.scala 48:55:@8411.4]
  wire [2:0] _T_9012; // @[Bitwise.scala 48:55:@8412.4]
  wire [3:0] _T_9013; // @[Bitwise.scala 48:55:@8413.4]
  wire [4:0] _T_9014; // @[Bitwise.scala 48:55:@8414.4]
  wire [1:0] _T_9015; // @[Bitwise.scala 48:55:@8415.4]
  wire [1:0] _T_9016; // @[Bitwise.scala 48:55:@8416.4]
  wire [2:0] _T_9017; // @[Bitwise.scala 48:55:@8417.4]
  wire [1:0] _T_9018; // @[Bitwise.scala 48:55:@8418.4]
  wire [1:0] _T_9019; // @[Bitwise.scala 48:55:@8419.4]
  wire [2:0] _T_9020; // @[Bitwise.scala 48:55:@8420.4]
  wire [3:0] _T_9021; // @[Bitwise.scala 48:55:@8421.4]
  wire [1:0] _T_9022; // @[Bitwise.scala 48:55:@8422.4]
  wire [1:0] _T_9023; // @[Bitwise.scala 48:55:@8423.4]
  wire [2:0] _T_9024; // @[Bitwise.scala 48:55:@8424.4]
  wire [1:0] _T_9025; // @[Bitwise.scala 48:55:@8425.4]
  wire [1:0] _T_9026; // @[Bitwise.scala 48:55:@8426.4]
  wire [2:0] _T_9027; // @[Bitwise.scala 48:55:@8427.4]
  wire [3:0] _T_9028; // @[Bitwise.scala 48:55:@8428.4]
  wire [4:0] _T_9029; // @[Bitwise.scala 48:55:@8429.4]
  wire [5:0] _T_9030; // @[Bitwise.scala 48:55:@8430.4]
  wire [1:0] _T_9031; // @[Bitwise.scala 48:55:@8431.4]
  wire [1:0] _T_9032; // @[Bitwise.scala 48:55:@8432.4]
  wire [2:0] _T_9033; // @[Bitwise.scala 48:55:@8433.4]
  wire [1:0] _T_9034; // @[Bitwise.scala 48:55:@8434.4]
  wire [1:0] _T_9035; // @[Bitwise.scala 48:55:@8435.4]
  wire [2:0] _T_9036; // @[Bitwise.scala 48:55:@8436.4]
  wire [3:0] _T_9037; // @[Bitwise.scala 48:55:@8437.4]
  wire [1:0] _T_9038; // @[Bitwise.scala 48:55:@8438.4]
  wire [1:0] _T_9039; // @[Bitwise.scala 48:55:@8439.4]
  wire [2:0] _T_9040; // @[Bitwise.scala 48:55:@8440.4]
  wire [1:0] _T_9041; // @[Bitwise.scala 48:55:@8441.4]
  wire [1:0] _T_9042; // @[Bitwise.scala 48:55:@8442.4]
  wire [2:0] _T_9043; // @[Bitwise.scala 48:55:@8443.4]
  wire [3:0] _T_9044; // @[Bitwise.scala 48:55:@8444.4]
  wire [4:0] _T_9045; // @[Bitwise.scala 48:55:@8445.4]
  wire [1:0] _T_9046; // @[Bitwise.scala 48:55:@8446.4]
  wire [1:0] _T_9047; // @[Bitwise.scala 48:55:@8447.4]
  wire [2:0] _T_9048; // @[Bitwise.scala 48:55:@8448.4]
  wire [1:0] _T_9049; // @[Bitwise.scala 48:55:@8449.4]
  wire [1:0] _T_9050; // @[Bitwise.scala 48:55:@8450.4]
  wire [2:0] _T_9051; // @[Bitwise.scala 48:55:@8451.4]
  wire [3:0] _T_9052; // @[Bitwise.scala 48:55:@8452.4]
  wire [1:0] _T_9053; // @[Bitwise.scala 48:55:@8453.4]
  wire [1:0] _T_9054; // @[Bitwise.scala 48:55:@8454.4]
  wire [2:0] _T_9055; // @[Bitwise.scala 48:55:@8455.4]
  wire [1:0] _T_9056; // @[Bitwise.scala 48:55:@8456.4]
  wire [1:0] _T_9057; // @[Bitwise.scala 48:55:@8457.4]
  wire [2:0] _T_9058; // @[Bitwise.scala 48:55:@8458.4]
  wire [3:0] _T_9059; // @[Bitwise.scala 48:55:@8459.4]
  wire [4:0] _T_9060; // @[Bitwise.scala 48:55:@8460.4]
  wire [5:0] _T_9061; // @[Bitwise.scala 48:55:@8461.4]
  wire [6:0] _T_9062; // @[Bitwise.scala 48:55:@8462.4]
  wire  _T_9128; // @[Bitwise.scala 50:65:@8529.4]
  wire  _T_9129; // @[Bitwise.scala 50:65:@8530.4]
  wire  _T_9130; // @[Bitwise.scala 50:65:@8531.4]
  wire  _T_9131; // @[Bitwise.scala 50:65:@8532.4]
  wire  _T_9132; // @[Bitwise.scala 50:65:@8533.4]
  wire  _T_9133; // @[Bitwise.scala 50:65:@8534.4]
  wire  _T_9134; // @[Bitwise.scala 50:65:@8535.4]
  wire  _T_9135; // @[Bitwise.scala 50:65:@8536.4]
  wire  _T_9136; // @[Bitwise.scala 50:65:@8537.4]
  wire  _T_9137; // @[Bitwise.scala 50:65:@8538.4]
  wire  _T_9138; // @[Bitwise.scala 50:65:@8539.4]
  wire  _T_9139; // @[Bitwise.scala 50:65:@8540.4]
  wire  _T_9140; // @[Bitwise.scala 50:65:@8541.4]
  wire  _T_9141; // @[Bitwise.scala 50:65:@8542.4]
  wire  _T_9142; // @[Bitwise.scala 50:65:@8543.4]
  wire  _T_9143; // @[Bitwise.scala 50:65:@8544.4]
  wire  _T_9144; // @[Bitwise.scala 50:65:@8545.4]
  wire  _T_9145; // @[Bitwise.scala 50:65:@8546.4]
  wire  _T_9146; // @[Bitwise.scala 50:65:@8547.4]
  wire  _T_9147; // @[Bitwise.scala 50:65:@8548.4]
  wire  _T_9148; // @[Bitwise.scala 50:65:@8549.4]
  wire  _T_9149; // @[Bitwise.scala 50:65:@8550.4]
  wire  _T_9150; // @[Bitwise.scala 50:65:@8551.4]
  wire  _T_9151; // @[Bitwise.scala 50:65:@8552.4]
  wire  _T_9152; // @[Bitwise.scala 50:65:@8553.4]
  wire  _T_9153; // @[Bitwise.scala 50:65:@8554.4]
  wire  _T_9154; // @[Bitwise.scala 50:65:@8555.4]
  wire  _T_9155; // @[Bitwise.scala 50:65:@8556.4]
  wire  _T_9156; // @[Bitwise.scala 50:65:@8557.4]
  wire  _T_9157; // @[Bitwise.scala 50:65:@8558.4]
  wire  _T_9158; // @[Bitwise.scala 50:65:@8559.4]
  wire  _T_9159; // @[Bitwise.scala 50:65:@8560.4]
  wire  _T_9160; // @[Bitwise.scala 50:65:@8561.4]
  wire  _T_9161; // @[Bitwise.scala 50:65:@8562.4]
  wire  _T_9162; // @[Bitwise.scala 50:65:@8563.4]
  wire  _T_9163; // @[Bitwise.scala 50:65:@8564.4]
  wire  _T_9164; // @[Bitwise.scala 50:65:@8565.4]
  wire  _T_9165; // @[Bitwise.scala 50:65:@8566.4]
  wire  _T_9166; // @[Bitwise.scala 50:65:@8567.4]
  wire  _T_9167; // @[Bitwise.scala 50:65:@8568.4]
  wire  _T_9168; // @[Bitwise.scala 50:65:@8569.4]
  wire  _T_9169; // @[Bitwise.scala 50:65:@8570.4]
  wire  _T_9170; // @[Bitwise.scala 50:65:@8571.4]
  wire  _T_9171; // @[Bitwise.scala 50:65:@8572.4]
  wire  _T_9172; // @[Bitwise.scala 50:65:@8573.4]
  wire  _T_9173; // @[Bitwise.scala 50:65:@8574.4]
  wire  _T_9174; // @[Bitwise.scala 50:65:@8575.4]
  wire  _T_9175; // @[Bitwise.scala 50:65:@8576.4]
  wire  _T_9176; // @[Bitwise.scala 50:65:@8577.4]
  wire  _T_9177; // @[Bitwise.scala 50:65:@8578.4]
  wire  _T_9178; // @[Bitwise.scala 50:65:@8579.4]
  wire  _T_9179; // @[Bitwise.scala 50:65:@8580.4]
  wire  _T_9180; // @[Bitwise.scala 50:65:@8581.4]
  wire  _T_9181; // @[Bitwise.scala 50:65:@8582.4]
  wire  _T_9182; // @[Bitwise.scala 50:65:@8583.4]
  wire  _T_9183; // @[Bitwise.scala 50:65:@8584.4]
  wire  _T_9184; // @[Bitwise.scala 50:65:@8585.4]
  wire  _T_9185; // @[Bitwise.scala 50:65:@8586.4]
  wire  _T_9186; // @[Bitwise.scala 50:65:@8587.4]
  wire  _T_9187; // @[Bitwise.scala 50:65:@8588.4]
  wire  _T_9188; // @[Bitwise.scala 50:65:@8589.4]
  wire  _T_9189; // @[Bitwise.scala 50:65:@8590.4]
  wire  _T_9190; // @[Bitwise.scala 50:65:@8591.4]
  wire [1:0] _T_9191; // @[Bitwise.scala 48:55:@8592.4]
  wire [1:0] _T_9192; // @[Bitwise.scala 48:55:@8593.4]
  wire [2:0] _T_9193; // @[Bitwise.scala 48:55:@8594.4]
  wire [1:0] _T_9194; // @[Bitwise.scala 48:55:@8595.4]
  wire [1:0] _T_9195; // @[Bitwise.scala 48:55:@8596.4]
  wire [2:0] _T_9196; // @[Bitwise.scala 48:55:@8597.4]
  wire [3:0] _T_9197; // @[Bitwise.scala 48:55:@8598.4]
  wire [1:0] _T_9198; // @[Bitwise.scala 48:55:@8599.4]
  wire [1:0] _T_9199; // @[Bitwise.scala 48:55:@8600.4]
  wire [2:0] _T_9200; // @[Bitwise.scala 48:55:@8601.4]
  wire [1:0] _T_9201; // @[Bitwise.scala 48:55:@8602.4]
  wire [1:0] _T_9202; // @[Bitwise.scala 48:55:@8603.4]
  wire [2:0] _T_9203; // @[Bitwise.scala 48:55:@8604.4]
  wire [3:0] _T_9204; // @[Bitwise.scala 48:55:@8605.4]
  wire [4:0] _T_9205; // @[Bitwise.scala 48:55:@8606.4]
  wire [1:0] _T_9206; // @[Bitwise.scala 48:55:@8607.4]
  wire [1:0] _T_9207; // @[Bitwise.scala 48:55:@8608.4]
  wire [2:0] _T_9208; // @[Bitwise.scala 48:55:@8609.4]
  wire [1:0] _T_9209; // @[Bitwise.scala 48:55:@8610.4]
  wire [1:0] _T_9210; // @[Bitwise.scala 48:55:@8611.4]
  wire [2:0] _T_9211; // @[Bitwise.scala 48:55:@8612.4]
  wire [3:0] _T_9212; // @[Bitwise.scala 48:55:@8613.4]
  wire [1:0] _T_9213; // @[Bitwise.scala 48:55:@8614.4]
  wire [1:0] _T_9214; // @[Bitwise.scala 48:55:@8615.4]
  wire [2:0] _T_9215; // @[Bitwise.scala 48:55:@8616.4]
  wire [1:0] _T_9216; // @[Bitwise.scala 48:55:@8617.4]
  wire [1:0] _T_9217; // @[Bitwise.scala 48:55:@8618.4]
  wire [2:0] _T_9218; // @[Bitwise.scala 48:55:@8619.4]
  wire [3:0] _T_9219; // @[Bitwise.scala 48:55:@8620.4]
  wire [4:0] _T_9220; // @[Bitwise.scala 48:55:@8621.4]
  wire [5:0] _T_9221; // @[Bitwise.scala 48:55:@8622.4]
  wire [1:0] _T_9222; // @[Bitwise.scala 48:55:@8623.4]
  wire [1:0] _T_9223; // @[Bitwise.scala 48:55:@8624.4]
  wire [2:0] _T_9224; // @[Bitwise.scala 48:55:@8625.4]
  wire [1:0] _T_9225; // @[Bitwise.scala 48:55:@8626.4]
  wire [1:0] _T_9226; // @[Bitwise.scala 48:55:@8627.4]
  wire [2:0] _T_9227; // @[Bitwise.scala 48:55:@8628.4]
  wire [3:0] _T_9228; // @[Bitwise.scala 48:55:@8629.4]
  wire [1:0] _T_9229; // @[Bitwise.scala 48:55:@8630.4]
  wire [1:0] _T_9230; // @[Bitwise.scala 48:55:@8631.4]
  wire [2:0] _T_9231; // @[Bitwise.scala 48:55:@8632.4]
  wire [1:0] _T_9232; // @[Bitwise.scala 48:55:@8633.4]
  wire [1:0] _T_9233; // @[Bitwise.scala 48:55:@8634.4]
  wire [2:0] _T_9234; // @[Bitwise.scala 48:55:@8635.4]
  wire [3:0] _T_9235; // @[Bitwise.scala 48:55:@8636.4]
  wire [4:0] _T_9236; // @[Bitwise.scala 48:55:@8637.4]
  wire [1:0] _T_9237; // @[Bitwise.scala 48:55:@8638.4]
  wire [1:0] _T_9238; // @[Bitwise.scala 48:55:@8639.4]
  wire [2:0] _T_9239; // @[Bitwise.scala 48:55:@8640.4]
  wire [1:0] _T_9240; // @[Bitwise.scala 48:55:@8641.4]
  wire [1:0] _T_9241; // @[Bitwise.scala 48:55:@8642.4]
  wire [2:0] _T_9242; // @[Bitwise.scala 48:55:@8643.4]
  wire [3:0] _T_9243; // @[Bitwise.scala 48:55:@8644.4]
  wire [1:0] _T_9244; // @[Bitwise.scala 48:55:@8645.4]
  wire [1:0] _T_9245; // @[Bitwise.scala 48:55:@8646.4]
  wire [2:0] _T_9246; // @[Bitwise.scala 48:55:@8647.4]
  wire [1:0] _T_9247; // @[Bitwise.scala 48:55:@8648.4]
  wire [1:0] _T_9248; // @[Bitwise.scala 48:55:@8649.4]
  wire [2:0] _T_9249; // @[Bitwise.scala 48:55:@8650.4]
  wire [3:0] _T_9250; // @[Bitwise.scala 48:55:@8651.4]
  wire [4:0] _T_9251; // @[Bitwise.scala 48:55:@8652.4]
  wire [5:0] _T_9252; // @[Bitwise.scala 48:55:@8653.4]
  wire [6:0] _T_9253; // @[Bitwise.scala 48:55:@8654.4]
  reg  _T_9256; // @[NV_NVDLA_CSC_WL_dec.scala 89:27:@8656.4]
  reg [31:0] _RAND_0;
  reg [7:0] _T_9260_0; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_1;
  reg [7:0] _T_9260_1; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_2;
  reg [7:0] _T_9260_2; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_9260_3; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_4;
  reg [7:0] _T_9260_4; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_5;
  reg [7:0] _T_9260_5; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_6;
  reg [7:0] _T_9260_6; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_7;
  reg [7:0] _T_9260_7; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_9260_8; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_9260_9; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_10;
  reg [7:0] _T_9260_10; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_9260_11; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_9260_12; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_13;
  reg [7:0] _T_9260_13; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_14;
  reg [7:0] _T_9260_14; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_15;
  reg [7:0] _T_9260_15; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_16;
  reg [7:0] _T_9260_16; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_17;
  reg [7:0] _T_9260_17; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_18;
  reg [7:0] _T_9260_18; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_19;
  reg [7:0] _T_9260_19; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_9260_20; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_9260_21; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_9260_22; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_9260_23; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_9260_24; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_9260_25; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_9260_26; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_9260_27; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_28;
  reg [7:0] _T_9260_28; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_9260_29; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_9260_30; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_9260_31; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_9260_32; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_33;
  reg [7:0] _T_9260_33; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_9260_34; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_9260_35; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_9260_36; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_9260_37; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_38;
  reg [7:0] _T_9260_38; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_9260_39; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_9260_40; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_9260_41; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_9260_42; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_43;
  reg [7:0] _T_9260_43; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_9260_44; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_9260_45; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_9260_46; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_9260_47; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_48;
  reg [7:0] _T_9260_48; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_49;
  reg [7:0] _T_9260_49; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_50;
  reg [7:0] _T_9260_50; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_51;
  reg [7:0] _T_9260_51; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_52;
  reg [7:0] _T_9260_52; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_53;
  reg [7:0] _T_9260_53; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_9260_54; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_55;
  reg [7:0] _T_9260_55; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_56;
  reg [7:0] _T_9260_56; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_57;
  reg [7:0] _T_9260_57; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_58;
  reg [7:0] _T_9260_58; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_59;
  reg [7:0] _T_9260_59; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_9260_60; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_61;
  reg [7:0] _T_9260_61; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_62;
  reg [7:0] _T_9260_62; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_63;
  reg [7:0] _T_9260_63; // @[NV_NVDLA_CSC_WL_dec.scala 90:22:@8657.4]
  reg [31:0] _RAND_64;
  reg  _T_9330_0; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_65;
  reg  _T_9330_1; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_66;
  reg  _T_9330_2; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_67;
  reg  _T_9330_3; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_68;
  reg  _T_9330_4; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_69;
  reg  _T_9330_5; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_70;
  reg  _T_9330_6; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_71;
  reg  _T_9330_7; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_72;
  reg  _T_9330_8; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_73;
  reg  _T_9330_9; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_74;
  reg  _T_9330_10; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_75;
  reg  _T_9330_11; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_76;
  reg  _T_9330_12; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_77;
  reg  _T_9330_13; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_78;
  reg  _T_9330_14; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_79;
  reg  _T_9330_15; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_80;
  reg  _T_9330_16; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_81;
  reg  _T_9330_17; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_82;
  reg  _T_9330_18; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_83;
  reg  _T_9330_19; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_84;
  reg  _T_9330_20; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_85;
  reg  _T_9330_21; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_86;
  reg  _T_9330_22; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_87;
  reg  _T_9330_23; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_88;
  reg  _T_9330_24; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_89;
  reg  _T_9330_25; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_90;
  reg  _T_9330_26; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_91;
  reg  _T_9330_27; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_92;
  reg  _T_9330_28; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_93;
  reg  _T_9330_29; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_94;
  reg  _T_9330_30; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_95;
  reg  _T_9330_31; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_96;
  reg  _T_9330_32; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_97;
  reg  _T_9330_33; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_98;
  reg  _T_9330_34; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_99;
  reg  _T_9330_35; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_100;
  reg  _T_9330_36; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_101;
  reg  _T_9330_37; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_102;
  reg  _T_9330_38; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_103;
  reg  _T_9330_39; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_104;
  reg  _T_9330_40; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_105;
  reg  _T_9330_41; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_106;
  reg  _T_9330_42; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_107;
  reg  _T_9330_43; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_108;
  reg  _T_9330_44; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_109;
  reg  _T_9330_45; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_110;
  reg  _T_9330_46; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_111;
  reg  _T_9330_47; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_112;
  reg  _T_9330_48; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_113;
  reg  _T_9330_49; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_114;
  reg  _T_9330_50; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_115;
  reg  _T_9330_51; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_116;
  reg  _T_9330_52; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_117;
  reg  _T_9330_53; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_118;
  reg  _T_9330_54; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_119;
  reg  _T_9330_55; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_120;
  reg  _T_9330_56; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_121;
  reg  _T_9330_57; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_122;
  reg  _T_9330_58; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_123;
  reg  _T_9330_59; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_124;
  reg  _T_9330_60; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_125;
  reg  _T_9330_61; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_126;
  reg  _T_9330_62; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_127;
  reg  _T_9330_63; // @[NV_NVDLA_CSC_WL_dec.scala 91:22:@8658.4]
  reg [31:0] _RAND_128;
  reg  _T_9535_0; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_129;
  reg  _T_9535_1; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_130;
  reg  _T_9535_2; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_131;
  reg  _T_9535_3; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_132;
  reg  _T_9535_4; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_133;
  reg  _T_9535_5; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_134;
  reg  _T_9535_6; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_135;
  reg  _T_9535_7; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_136;
  reg  _T_9535_8; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_137;
  reg  _T_9535_9; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_138;
  reg  _T_9535_10; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_139;
  reg  _T_9535_11; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_140;
  reg  _T_9535_12; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_141;
  reg  _T_9535_13; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_142;
  reg  _T_9535_14; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_143;
  reg  _T_9535_15; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_144;
  reg  _T_9535_16; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_145;
  reg  _T_9535_17; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_146;
  reg  _T_9535_18; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_147;
  reg  _T_9535_19; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_148;
  reg  _T_9535_20; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_149;
  reg  _T_9535_21; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_150;
  reg  _T_9535_22; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_151;
  reg  _T_9535_23; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_152;
  reg  _T_9535_24; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_153;
  reg  _T_9535_25; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_154;
  reg  _T_9535_26; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_155;
  reg  _T_9535_27; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_156;
  reg  _T_9535_28; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_157;
  reg  _T_9535_29; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_158;
  reg  _T_9535_30; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_159;
  reg  _T_9535_31; // @[NV_NVDLA_CSC_WL_dec.scala 92:25:@8692.4]
  reg [31:0] _RAND_160;
  reg [6:0] _T_10211_63; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_161;
  reg [5:0] _T_10211_62; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_162;
  reg [5:0] _T_10211_61; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_163;
  reg [5:0] _T_10211_60; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_164;
  reg [5:0] _T_10211_59; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_165;
  reg [5:0] _T_10211_58; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_166;
  reg [5:0] _T_10211_57; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_167;
  reg [5:0] _T_10211_56; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_168;
  reg [5:0] _T_10211_55; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_169;
  reg [5:0] _T_10211_54; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_170;
  reg [5:0] _T_10211_53; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_171;
  reg [5:0] _T_10211_52; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_172;
  reg [5:0] _T_10211_51; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_173;
  reg [5:0] _T_10211_50; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_174;
  reg [5:0] _T_10211_49; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_175;
  reg [5:0] _T_10211_48; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_176;
  reg [5:0] _T_10211_47; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_177;
  reg [5:0] _T_10211_46; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_178;
  reg [5:0] _T_10211_45; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_179;
  reg [5:0] _T_10211_44; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_180;
  reg [5:0] _T_10211_43; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_181;
  reg [5:0] _T_10211_42; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_182;
  reg [5:0] _T_10211_41; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_183;
  reg [5:0] _T_10211_40; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_184;
  reg [5:0] _T_10211_39; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_185;
  reg [5:0] _T_10211_38; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_186;
  reg [5:0] _T_10211_37; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_187;
  reg [5:0] _T_10211_36; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_188;
  reg [5:0] _T_10211_35; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_189;
  reg [5:0] _T_10211_34; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_190;
  reg [5:0] _T_10211_33; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_191;
  reg [5:0] _T_10211_32; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_192;
  reg [5:0] _T_10211_31; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_193;
  reg [4:0] _T_10211_30; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_194;
  reg [4:0] _T_10211_29; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_195;
  reg [4:0] _T_10211_28; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_196;
  reg [4:0] _T_10211_27; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_197;
  reg [4:0] _T_10211_26; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_198;
  reg [4:0] _T_10211_25; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_199;
  reg [4:0] _T_10211_24; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_200;
  reg [4:0] _T_10211_23; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_201;
  reg [4:0] _T_10211_22; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_202;
  reg [4:0] _T_10211_21; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_203;
  reg [4:0] _T_10211_20; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_204;
  reg [4:0] _T_10211_19; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_205;
  reg [4:0] _T_10211_18; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_206;
  reg [4:0] _T_10211_17; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_207;
  reg [4:0] _T_10211_16; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_208;
  reg [4:0] _T_10211_15; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_209;
  reg [3:0] _T_10211_14; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_210;
  reg [3:0] _T_10211_13; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_211;
  reg [3:0] _T_10211_12; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_212;
  reg [3:0] _T_10211_11; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_213;
  reg [3:0] _T_10211_10; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_214;
  reg [3:0] _T_10211_9; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_215;
  reg [3:0] _T_10211_8; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_216;
  reg [3:0] _T_10211_7; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_217;
  reg [2:0] _T_10211_6; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_218;
  reg [2:0] _T_10211_5; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_219;
  reg [2:0] _T_10211_4; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_220;
  reg [2:0] _T_10211_3; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_221;
  reg [1:0] _T_10211_2; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_222;
  reg [1:0] _T_10211_1; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_223;
  reg  _T_10211_0; // @[NV_NVDLA_CSC_WL_dec.scala 93:29:@8821.4]
  reg [31:0] _RAND_224;
  wire  _GEN_128; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_129; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_130; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_131; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_132; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_133; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_134; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_135; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_136; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_137; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_138; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_139; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_140; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_141; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_142; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_143; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_144; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_145; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_146; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_147; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_148; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_149; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_150; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_151; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_152; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_153; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_154; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_155; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_156; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  wire  _T_10212; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@8985.4]
  wire  _T_10213; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@8986.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@8987.4]
  wire [1:0] _GEN_161; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@8992.4]
  wire [1:0] _T_1061_2; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@603.4]
  wire [1:0] _GEN_162; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@8997.4]
  wire [2:0] _GEN_163; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9002.4]
  wire [2:0] _T_1061_4; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@749.4]
  wire [2:0] _GEN_164; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9007.4]
  wire [2:0] _T_1061_5; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@825.4]
  wire [2:0] _GEN_165; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9012.4]
  wire [2:0] _T_1061_6; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@903.4]
  wire [2:0] _GEN_166; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9017.4]
  wire [3:0] _GEN_167; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9022.4]
  wire  _T_10228; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9025.4]
  wire  _T_10229; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9026.4]
  wire [3:0] _T_1061_8; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1065.4]
  wire [3:0] _GEN_168; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9027.4]
  wire [3:0] _T_1061_9; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1149.4]
  wire [3:0] _GEN_169; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9032.4]
  wire [3:0] _T_1061_10; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1235.4]
  wire [3:0] _GEN_170; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9037.4]
  wire [3:0] _T_1061_11; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1323.4]
  wire [3:0] _GEN_171; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9042.4]
  wire [3:0] _T_1061_12; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1413.4]
  wire [3:0] _GEN_172; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9047.4]
  wire [3:0] _T_1061_13; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1505.4]
  wire [3:0] _GEN_173; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9052.4]
  wire [3:0] _T_1061_14; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1599.4]
  wire [3:0] _GEN_174; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9057.4]
  wire [4:0] _GEN_175; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9062.4]
  wire  _T_10244; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9065.4]
  wire  _T_10245; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9066.4]
  wire [4:0] _T_1061_16; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1793.4]
  wire [4:0] _GEN_176; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9067.4]
  wire [4:0] _T_1061_17; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1893.4]
  wire [4:0] _GEN_177; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9072.4]
  wire [4:0] _T_1061_18; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1995.4]
  wire [4:0] _GEN_178; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9077.4]
  wire [4:0] _T_1061_19; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2099.4]
  wire [4:0] _GEN_179; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9082.4]
  wire [4:0] _T_1061_20; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2205.4]
  wire [4:0] _GEN_180; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9087.4]
  wire [4:0] _T_1061_21; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2313.4]
  wire [4:0] _GEN_181; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9092.4]
  wire [4:0] _T_1061_22; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2423.4]
  wire [4:0] _GEN_182; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9097.4]
  wire [4:0] _T_1061_23; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2535.4]
  wire [4:0] _GEN_183; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9102.4]
  wire  _T_10260; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9105.4]
  wire  _T_10261; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9106.4]
  wire [4:0] _T_1061_24; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2649.4]
  wire [4:0] _GEN_184; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9107.4]
  wire [4:0] _T_1061_25; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2765.4]
  wire [4:0] _GEN_185; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9112.4]
  wire [4:0] _T_1061_26; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2883.4]
  wire [4:0] _GEN_186; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9117.4]
  wire [4:0] _T_1061_27; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3003.4]
  wire [4:0] _GEN_187; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9122.4]
  wire [4:0] _T_1061_28; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3125.4]
  wire [4:0] _GEN_188; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9127.4]
  wire [4:0] _T_1061_29; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3249.4]
  wire [4:0] _GEN_189; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9132.4]
  wire [4:0] _T_1061_30; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3375.4]
  wire [4:0] _GEN_190; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9137.4]
  wire [5:0] _GEN_191; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9142.4]
  wire  _T_10276; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9145.4]
  wire  _T_10277; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9146.4]
  wire [5:0] _T_1061_32; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3633.4]
  wire [5:0] _GEN_192; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9147.4]
  wire [5:0] _T_1061_33; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3765.4]
  wire [5:0] _GEN_193; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9152.4]
  wire [5:0] _T_1061_34; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3899.4]
  wire [5:0] _GEN_194; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9157.4]
  wire [5:0] _T_1061_35; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4035.4]
  wire [5:0] _GEN_195; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9162.4]
  wire [5:0] _T_1061_36; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4173.4]
  wire [5:0] _GEN_196; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9167.4]
  wire [5:0] _T_1061_37; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4313.4]
  wire [5:0] _GEN_197; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9172.4]
  wire [5:0] _T_1061_38; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4455.4]
  wire [5:0] _GEN_198; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9177.4]
  wire [5:0] _T_1061_39; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4599.4]
  wire [5:0] _GEN_199; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9182.4]
  wire  _T_10292; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9185.4]
  wire  _T_10293; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9186.4]
  wire [5:0] _T_1061_40; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4745.4]
  wire [5:0] _GEN_200; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9187.4]
  wire [5:0] _T_1061_41; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4893.4]
  wire [5:0] _GEN_201; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9192.4]
  wire [5:0] _T_1061_42; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5043.4]
  wire [5:0] _GEN_202; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9197.4]
  wire [5:0] _T_1061_43; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5195.4]
  wire [5:0] _GEN_203; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9202.4]
  wire [5:0] _T_1061_44; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5349.4]
  wire [5:0] _GEN_204; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9207.4]
  wire [5:0] _T_1061_45; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5505.4]
  wire [5:0] _GEN_205; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9212.4]
  wire [5:0] _T_1061_46; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5663.4]
  wire [5:0] _GEN_206; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9217.4]
  wire [5:0] _T_1061_47; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5823.4]
  wire [5:0] _GEN_207; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9222.4]
  wire  _T_10308; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9225.4]
  wire  _T_10309; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9226.4]
  wire [5:0] _T_1061_48; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5985.4]
  wire [5:0] _GEN_208; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9227.4]
  wire [5:0] _T_1061_49; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6149.4]
  wire [5:0] _GEN_209; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9232.4]
  wire [5:0] _T_1061_50; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6315.4]
  wire [5:0] _GEN_210; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9237.4]
  wire [5:0] _T_1061_51; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6483.4]
  wire [5:0] _GEN_211; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9242.4]
  wire [5:0] _T_1061_52; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6653.4]
  wire [5:0] _GEN_212; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9247.4]
  wire [5:0] _T_1061_53; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6825.4]
  wire [5:0] _GEN_213; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9252.4]
  wire [5:0] _T_1061_54; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6999.4]
  wire [5:0] _GEN_214; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9257.4]
  wire [5:0] _T_1061_55; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7175.4]
  wire [5:0] _GEN_215; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9262.4]
  wire  _T_10324; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9265.4]
  wire  _T_10325; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9266.4]
  wire [5:0] _T_1061_56; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7353.4]
  wire [5:0] _GEN_216; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9267.4]
  wire [5:0] _T_1061_57; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7533.4]
  wire [5:0] _GEN_217; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9272.4]
  wire [5:0] _T_1061_58; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7715.4]
  wire [5:0] _GEN_218; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9277.4]
  wire [5:0] _T_1061_59; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7899.4]
  wire [5:0] _GEN_219; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9282.4]
  wire [5:0] _T_1061_60; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@8085.4]
  wire [5:0] _GEN_220; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9287.4]
  wire [5:0] _T_1061_61; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@8273.4]
  wire [5:0] _GEN_221; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9292.4]
  wire [5:0] _T_1061_62; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@8463.4]
  wire [5:0] _GEN_222; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9297.4]
  wire [6:0] _GEN_223; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9302.4]
  wire [7:0] _T_10413; // @[Mux.scala 46:16:@9307.4]
  wire  _T_10417; // @[Mux.scala 46:19:@9309.4]
  wire [7:0] _T_10418; // @[Mux.scala 46:16:@9310.4]
  wire  _T_10419; // @[Mux.scala 46:19:@9311.4]
  wire [7:0] _T_10420; // @[Mux.scala 46:16:@9312.4]
  wire  _T_10425; // @[Mux.scala 46:19:@9314.4]
  wire [7:0] _T_10426; // @[Mux.scala 46:16:@9315.4]
  wire  _T_10427; // @[Mux.scala 46:19:@9316.4]
  wire [7:0] _T_10428; // @[Mux.scala 46:16:@9317.4]
  wire  _T_10429; // @[Mux.scala 46:19:@9318.4]
  wire [7:0] _T_10430; // @[Mux.scala 46:16:@9319.4]
  wire  _T_10436; // @[Mux.scala 46:19:@9321.4]
  wire [7:0] _T_10437; // @[Mux.scala 46:16:@9322.4]
  wire  _T_10438; // @[Mux.scala 46:19:@9323.4]
  wire [7:0] _T_10439; // @[Mux.scala 46:16:@9324.4]
  wire  _T_10440; // @[Mux.scala 46:19:@9325.4]
  wire [7:0] _T_10441; // @[Mux.scala 46:16:@9326.4]
  wire  _T_10442; // @[Mux.scala 46:19:@9327.4]
  wire [7:0] _T_10443; // @[Mux.scala 46:16:@9328.4]
  wire  _T_10450; // @[Mux.scala 46:19:@9330.4]
  wire [7:0] _T_10451; // @[Mux.scala 46:16:@9331.4]
  wire  _T_10452; // @[Mux.scala 46:19:@9332.4]
  wire [7:0] _T_10453; // @[Mux.scala 46:16:@9333.4]
  wire  _T_10454; // @[Mux.scala 46:19:@9334.4]
  wire [7:0] _T_10455; // @[Mux.scala 46:16:@9335.4]
  wire  _T_10456; // @[Mux.scala 46:19:@9336.4]
  wire [7:0] _T_10457; // @[Mux.scala 46:16:@9337.4]
  wire  _T_10458; // @[Mux.scala 46:19:@9338.4]
  wire [7:0] _T_10459; // @[Mux.scala 46:16:@9339.4]
  wire  _T_10467; // @[Mux.scala 46:19:@9341.4]
  wire [7:0] _T_10468; // @[Mux.scala 46:16:@9342.4]
  wire  _T_10469; // @[Mux.scala 46:19:@9343.4]
  wire [7:0] _T_10470; // @[Mux.scala 46:16:@9344.4]
  wire  _T_10471; // @[Mux.scala 46:19:@9345.4]
  wire [7:0] _T_10472; // @[Mux.scala 46:16:@9346.4]
  wire  _T_10473; // @[Mux.scala 46:19:@9347.4]
  wire [7:0] _T_10474; // @[Mux.scala 46:16:@9348.4]
  wire  _T_10475; // @[Mux.scala 46:19:@9349.4]
  wire [7:0] _T_10476; // @[Mux.scala 46:16:@9350.4]
  wire  _T_10477; // @[Mux.scala 46:19:@9351.4]
  wire [7:0] _T_10478; // @[Mux.scala 46:16:@9352.4]
  wire  _T_10487; // @[Mux.scala 46:19:@9354.4]
  wire [7:0] _T_10488; // @[Mux.scala 46:16:@9355.4]
  wire  _T_10489; // @[Mux.scala 46:19:@9356.4]
  wire [7:0] _T_10490; // @[Mux.scala 46:16:@9357.4]
  wire  _T_10491; // @[Mux.scala 46:19:@9358.4]
  wire [7:0] _T_10492; // @[Mux.scala 46:16:@9359.4]
  wire  _T_10493; // @[Mux.scala 46:19:@9360.4]
  wire [7:0] _T_10494; // @[Mux.scala 46:16:@9361.4]
  wire  _T_10495; // @[Mux.scala 46:19:@9362.4]
  wire [7:0] _T_10496; // @[Mux.scala 46:16:@9363.4]
  wire  _T_10497; // @[Mux.scala 46:19:@9364.4]
  wire [7:0] _T_10498; // @[Mux.scala 46:16:@9365.4]
  wire  _T_10499; // @[Mux.scala 46:19:@9366.4]
  wire [7:0] _T_10500; // @[Mux.scala 46:16:@9367.4]
  wire  _T_10510; // @[Mux.scala 46:19:@9369.4]
  wire [7:0] _T_10511; // @[Mux.scala 46:16:@9370.4]
  wire  _T_10512; // @[Mux.scala 46:19:@9371.4]
  wire [7:0] _T_10513; // @[Mux.scala 46:16:@9372.4]
  wire  _T_10514; // @[Mux.scala 46:19:@9373.4]
  wire [7:0] _T_10515; // @[Mux.scala 46:16:@9374.4]
  wire  _T_10516; // @[Mux.scala 46:19:@9375.4]
  wire [7:0] _T_10517; // @[Mux.scala 46:16:@9376.4]
  wire  _T_10518; // @[Mux.scala 46:19:@9377.4]
  wire [7:0] _T_10519; // @[Mux.scala 46:16:@9378.4]
  wire  _T_10520; // @[Mux.scala 46:19:@9379.4]
  wire [7:0] _T_10521; // @[Mux.scala 46:16:@9380.4]
  wire  _T_10522; // @[Mux.scala 46:19:@9381.4]
  wire [7:0] _T_10523; // @[Mux.scala 46:16:@9382.4]
  wire  _T_10524; // @[Mux.scala 46:19:@9383.4]
  wire [7:0] _T_10525; // @[Mux.scala 46:16:@9384.4]
  wire  _T_10536; // @[Mux.scala 46:19:@9386.4]
  wire [7:0] _T_10537; // @[Mux.scala 46:16:@9387.4]
  wire  _T_10538; // @[Mux.scala 46:19:@9388.4]
  wire [7:0] _T_10539; // @[Mux.scala 46:16:@9389.4]
  wire  _T_10540; // @[Mux.scala 46:19:@9390.4]
  wire [7:0] _T_10541; // @[Mux.scala 46:16:@9391.4]
  wire  _T_10542; // @[Mux.scala 46:19:@9392.4]
  wire [7:0] _T_10543; // @[Mux.scala 46:16:@9393.4]
  wire  _T_10544; // @[Mux.scala 46:19:@9394.4]
  wire [7:0] _T_10545; // @[Mux.scala 46:16:@9395.4]
  wire  _T_10546; // @[Mux.scala 46:19:@9396.4]
  wire [7:0] _T_10547; // @[Mux.scala 46:16:@9397.4]
  wire  _T_10548; // @[Mux.scala 46:19:@9398.4]
  wire [7:0] _T_10549; // @[Mux.scala 46:16:@9399.4]
  wire  _T_10550; // @[Mux.scala 46:19:@9400.4]
  wire [7:0] _T_10551; // @[Mux.scala 46:16:@9401.4]
  wire  _T_10552; // @[Mux.scala 46:19:@9402.4]
  wire [7:0] _T_10553; // @[Mux.scala 46:16:@9403.4]
  wire  _T_10565; // @[Mux.scala 46:19:@9405.4]
  wire [7:0] _T_10566; // @[Mux.scala 46:16:@9406.4]
  wire  _T_10567; // @[Mux.scala 46:19:@9407.4]
  wire [7:0] _T_10568; // @[Mux.scala 46:16:@9408.4]
  wire  _T_10569; // @[Mux.scala 46:19:@9409.4]
  wire [7:0] _T_10570; // @[Mux.scala 46:16:@9410.4]
  wire  _T_10571; // @[Mux.scala 46:19:@9411.4]
  wire [7:0] _T_10572; // @[Mux.scala 46:16:@9412.4]
  wire  _T_10573; // @[Mux.scala 46:19:@9413.4]
  wire [7:0] _T_10574; // @[Mux.scala 46:16:@9414.4]
  wire  _T_10575; // @[Mux.scala 46:19:@9415.4]
  wire [7:0] _T_10576; // @[Mux.scala 46:16:@9416.4]
  wire  _T_10577; // @[Mux.scala 46:19:@9417.4]
  wire [7:0] _T_10578; // @[Mux.scala 46:16:@9418.4]
  wire  _T_10579; // @[Mux.scala 46:19:@9419.4]
  wire [7:0] _T_10580; // @[Mux.scala 46:16:@9420.4]
  wire  _T_10581; // @[Mux.scala 46:19:@9421.4]
  wire [7:0] _T_10582; // @[Mux.scala 46:16:@9422.4]
  wire  _T_10583; // @[Mux.scala 46:19:@9423.4]
  wire [7:0] _T_10584; // @[Mux.scala 46:16:@9424.4]
  wire  _T_10597; // @[Mux.scala 46:19:@9426.4]
  wire [7:0] _T_10598; // @[Mux.scala 46:16:@9427.4]
  wire  _T_10599; // @[Mux.scala 46:19:@9428.4]
  wire [7:0] _T_10600; // @[Mux.scala 46:16:@9429.4]
  wire  _T_10601; // @[Mux.scala 46:19:@9430.4]
  wire [7:0] _T_10602; // @[Mux.scala 46:16:@9431.4]
  wire  _T_10603; // @[Mux.scala 46:19:@9432.4]
  wire [7:0] _T_10604; // @[Mux.scala 46:16:@9433.4]
  wire  _T_10605; // @[Mux.scala 46:19:@9434.4]
  wire [7:0] _T_10606; // @[Mux.scala 46:16:@9435.4]
  wire  _T_10607; // @[Mux.scala 46:19:@9436.4]
  wire [7:0] _T_10608; // @[Mux.scala 46:16:@9437.4]
  wire  _T_10609; // @[Mux.scala 46:19:@9438.4]
  wire [7:0] _T_10610; // @[Mux.scala 46:16:@9439.4]
  wire  _T_10611; // @[Mux.scala 46:19:@9440.4]
  wire [7:0] _T_10612; // @[Mux.scala 46:16:@9441.4]
  wire  _T_10613; // @[Mux.scala 46:19:@9442.4]
  wire [7:0] _T_10614; // @[Mux.scala 46:16:@9443.4]
  wire  _T_10615; // @[Mux.scala 46:19:@9444.4]
  wire [7:0] _T_10616; // @[Mux.scala 46:16:@9445.4]
  wire  _T_10617; // @[Mux.scala 46:19:@9446.4]
  wire [7:0] _T_10618; // @[Mux.scala 46:16:@9447.4]
  wire  _T_10632; // @[Mux.scala 46:19:@9449.4]
  wire [7:0] _T_10633; // @[Mux.scala 46:16:@9450.4]
  wire  _T_10634; // @[Mux.scala 46:19:@9451.4]
  wire [7:0] _T_10635; // @[Mux.scala 46:16:@9452.4]
  wire  _T_10636; // @[Mux.scala 46:19:@9453.4]
  wire [7:0] _T_10637; // @[Mux.scala 46:16:@9454.4]
  wire  _T_10638; // @[Mux.scala 46:19:@9455.4]
  wire [7:0] _T_10639; // @[Mux.scala 46:16:@9456.4]
  wire  _T_10640; // @[Mux.scala 46:19:@9457.4]
  wire [7:0] _T_10641; // @[Mux.scala 46:16:@9458.4]
  wire  _T_10642; // @[Mux.scala 46:19:@9459.4]
  wire [7:0] _T_10643; // @[Mux.scala 46:16:@9460.4]
  wire  _T_10644; // @[Mux.scala 46:19:@9461.4]
  wire [7:0] _T_10645; // @[Mux.scala 46:16:@9462.4]
  wire  _T_10646; // @[Mux.scala 46:19:@9463.4]
  wire [7:0] _T_10647; // @[Mux.scala 46:16:@9464.4]
  wire  _T_10648; // @[Mux.scala 46:19:@9465.4]
  wire [7:0] _T_10649; // @[Mux.scala 46:16:@9466.4]
  wire  _T_10650; // @[Mux.scala 46:19:@9467.4]
  wire [7:0] _T_10651; // @[Mux.scala 46:16:@9468.4]
  wire  _T_10652; // @[Mux.scala 46:19:@9469.4]
  wire [7:0] _T_10653; // @[Mux.scala 46:16:@9470.4]
  wire  _T_10654; // @[Mux.scala 46:19:@9471.4]
  wire [7:0] _T_10655; // @[Mux.scala 46:16:@9472.4]
  wire  _T_10670; // @[Mux.scala 46:19:@9474.4]
  wire [7:0] _T_10671; // @[Mux.scala 46:16:@9475.4]
  wire  _T_10672; // @[Mux.scala 46:19:@9476.4]
  wire [7:0] _T_10673; // @[Mux.scala 46:16:@9477.4]
  wire  _T_10674; // @[Mux.scala 46:19:@9478.4]
  wire [7:0] _T_10675; // @[Mux.scala 46:16:@9479.4]
  wire  _T_10676; // @[Mux.scala 46:19:@9480.4]
  wire [7:0] _T_10677; // @[Mux.scala 46:16:@9481.4]
  wire  _T_10678; // @[Mux.scala 46:19:@9482.4]
  wire [7:0] _T_10679; // @[Mux.scala 46:16:@9483.4]
  wire  _T_10680; // @[Mux.scala 46:19:@9484.4]
  wire [7:0] _T_10681; // @[Mux.scala 46:16:@9485.4]
  wire  _T_10682; // @[Mux.scala 46:19:@9486.4]
  wire [7:0] _T_10683; // @[Mux.scala 46:16:@9487.4]
  wire  _T_10684; // @[Mux.scala 46:19:@9488.4]
  wire [7:0] _T_10685; // @[Mux.scala 46:16:@9489.4]
  wire  _T_10686; // @[Mux.scala 46:19:@9490.4]
  wire [7:0] _T_10687; // @[Mux.scala 46:16:@9491.4]
  wire  _T_10688; // @[Mux.scala 46:19:@9492.4]
  wire [7:0] _T_10689; // @[Mux.scala 46:16:@9493.4]
  wire  _T_10690; // @[Mux.scala 46:19:@9494.4]
  wire [7:0] _T_10691; // @[Mux.scala 46:16:@9495.4]
  wire  _T_10692; // @[Mux.scala 46:19:@9496.4]
  wire [7:0] _T_10693; // @[Mux.scala 46:16:@9497.4]
  wire  _T_10694; // @[Mux.scala 46:19:@9498.4]
  wire [7:0] _T_10695; // @[Mux.scala 46:16:@9499.4]
  wire  _T_10711; // @[Mux.scala 46:19:@9501.4]
  wire [7:0] _T_10712; // @[Mux.scala 46:16:@9502.4]
  wire  _T_10713; // @[Mux.scala 46:19:@9503.4]
  wire [7:0] _T_10714; // @[Mux.scala 46:16:@9504.4]
  wire  _T_10715; // @[Mux.scala 46:19:@9505.4]
  wire [7:0] _T_10716; // @[Mux.scala 46:16:@9506.4]
  wire  _T_10717; // @[Mux.scala 46:19:@9507.4]
  wire [7:0] _T_10718; // @[Mux.scala 46:16:@9508.4]
  wire  _T_10719; // @[Mux.scala 46:19:@9509.4]
  wire [7:0] _T_10720; // @[Mux.scala 46:16:@9510.4]
  wire  _T_10721; // @[Mux.scala 46:19:@9511.4]
  wire [7:0] _T_10722; // @[Mux.scala 46:16:@9512.4]
  wire  _T_10723; // @[Mux.scala 46:19:@9513.4]
  wire [7:0] _T_10724; // @[Mux.scala 46:16:@9514.4]
  wire  _T_10725; // @[Mux.scala 46:19:@9515.4]
  wire [7:0] _T_10726; // @[Mux.scala 46:16:@9516.4]
  wire  _T_10727; // @[Mux.scala 46:19:@9517.4]
  wire [7:0] _T_10728; // @[Mux.scala 46:16:@9518.4]
  wire  _T_10729; // @[Mux.scala 46:19:@9519.4]
  wire [7:0] _T_10730; // @[Mux.scala 46:16:@9520.4]
  wire  _T_10731; // @[Mux.scala 46:19:@9521.4]
  wire [7:0] _T_10732; // @[Mux.scala 46:16:@9522.4]
  wire  _T_10733; // @[Mux.scala 46:19:@9523.4]
  wire [7:0] _T_10734; // @[Mux.scala 46:16:@9524.4]
  wire  _T_10735; // @[Mux.scala 46:19:@9525.4]
  wire [7:0] _T_10736; // @[Mux.scala 46:16:@9526.4]
  wire  _T_10737; // @[Mux.scala 46:19:@9527.4]
  wire [7:0] _T_10738; // @[Mux.scala 46:16:@9528.4]
  wire  _T_10755; // @[Mux.scala 46:19:@9530.4]
  wire [7:0] _T_10756; // @[Mux.scala 46:16:@9531.4]
  wire  _T_10757; // @[Mux.scala 46:19:@9532.4]
  wire [7:0] _T_10758; // @[Mux.scala 46:16:@9533.4]
  wire  _T_10759; // @[Mux.scala 46:19:@9534.4]
  wire [7:0] _T_10760; // @[Mux.scala 46:16:@9535.4]
  wire  _T_10761; // @[Mux.scala 46:19:@9536.4]
  wire [7:0] _T_10762; // @[Mux.scala 46:16:@9537.4]
  wire  _T_10763; // @[Mux.scala 46:19:@9538.4]
  wire [7:0] _T_10764; // @[Mux.scala 46:16:@9539.4]
  wire  _T_10765; // @[Mux.scala 46:19:@9540.4]
  wire [7:0] _T_10766; // @[Mux.scala 46:16:@9541.4]
  wire  _T_10767; // @[Mux.scala 46:19:@9542.4]
  wire [7:0] _T_10768; // @[Mux.scala 46:16:@9543.4]
  wire  _T_10769; // @[Mux.scala 46:19:@9544.4]
  wire [7:0] _T_10770; // @[Mux.scala 46:16:@9545.4]
  wire  _T_10771; // @[Mux.scala 46:19:@9546.4]
  wire [7:0] _T_10772; // @[Mux.scala 46:16:@9547.4]
  wire  _T_10773; // @[Mux.scala 46:19:@9548.4]
  wire [7:0] _T_10774; // @[Mux.scala 46:16:@9549.4]
  wire  _T_10775; // @[Mux.scala 46:19:@9550.4]
  wire [7:0] _T_10776; // @[Mux.scala 46:16:@9551.4]
  wire  _T_10777; // @[Mux.scala 46:19:@9552.4]
  wire [7:0] _T_10778; // @[Mux.scala 46:16:@9553.4]
  wire  _T_10779; // @[Mux.scala 46:19:@9554.4]
  wire [7:0] _T_10780; // @[Mux.scala 46:16:@9555.4]
  wire  _T_10781; // @[Mux.scala 46:19:@9556.4]
  wire [7:0] _T_10782; // @[Mux.scala 46:16:@9557.4]
  wire  _T_10783; // @[Mux.scala 46:19:@9558.4]
  wire [7:0] _T_10784; // @[Mux.scala 46:16:@9559.4]
  wire  _T_10802; // @[Mux.scala 46:19:@9561.4]
  wire [7:0] _T_10803; // @[Mux.scala 46:16:@9562.4]
  wire  _T_10804; // @[Mux.scala 46:19:@9563.4]
  wire [7:0] _T_10805; // @[Mux.scala 46:16:@9564.4]
  wire  _T_10806; // @[Mux.scala 46:19:@9565.4]
  wire [7:0] _T_10807; // @[Mux.scala 46:16:@9566.4]
  wire  _T_10808; // @[Mux.scala 46:19:@9567.4]
  wire [7:0] _T_10809; // @[Mux.scala 46:16:@9568.4]
  wire  _T_10810; // @[Mux.scala 46:19:@9569.4]
  wire [7:0] _T_10811; // @[Mux.scala 46:16:@9570.4]
  wire  _T_10812; // @[Mux.scala 46:19:@9571.4]
  wire [7:0] _T_10813; // @[Mux.scala 46:16:@9572.4]
  wire  _T_10814; // @[Mux.scala 46:19:@9573.4]
  wire [7:0] _T_10815; // @[Mux.scala 46:16:@9574.4]
  wire  _T_10816; // @[Mux.scala 46:19:@9575.4]
  wire [7:0] _T_10817; // @[Mux.scala 46:16:@9576.4]
  wire  _T_10818; // @[Mux.scala 46:19:@9577.4]
  wire [7:0] _T_10819; // @[Mux.scala 46:16:@9578.4]
  wire  _T_10820; // @[Mux.scala 46:19:@9579.4]
  wire [7:0] _T_10821; // @[Mux.scala 46:16:@9580.4]
  wire  _T_10822; // @[Mux.scala 46:19:@9581.4]
  wire [7:0] _T_10823; // @[Mux.scala 46:16:@9582.4]
  wire  _T_10824; // @[Mux.scala 46:19:@9583.4]
  wire [7:0] _T_10825; // @[Mux.scala 46:16:@9584.4]
  wire  _T_10826; // @[Mux.scala 46:19:@9585.4]
  wire [7:0] _T_10827; // @[Mux.scala 46:16:@9586.4]
  wire  _T_10828; // @[Mux.scala 46:19:@9587.4]
  wire [7:0] _T_10829; // @[Mux.scala 46:16:@9588.4]
  wire  _T_10830; // @[Mux.scala 46:19:@9589.4]
  wire [7:0] _T_10831; // @[Mux.scala 46:16:@9590.4]
  wire  _T_10832; // @[Mux.scala 46:19:@9591.4]
  wire [7:0] _T_10833; // @[Mux.scala 46:16:@9592.4]
  wire  _T_10852; // @[Mux.scala 46:19:@9594.4]
  wire [7:0] _T_10853; // @[Mux.scala 46:16:@9595.4]
  wire  _T_10854; // @[Mux.scala 46:19:@9596.4]
  wire [7:0] _T_10855; // @[Mux.scala 46:16:@9597.4]
  wire  _T_10856; // @[Mux.scala 46:19:@9598.4]
  wire [7:0] _T_10857; // @[Mux.scala 46:16:@9599.4]
  wire  _T_10858; // @[Mux.scala 46:19:@9600.4]
  wire [7:0] _T_10859; // @[Mux.scala 46:16:@9601.4]
  wire  _T_10860; // @[Mux.scala 46:19:@9602.4]
  wire [7:0] _T_10861; // @[Mux.scala 46:16:@9603.4]
  wire  _T_10862; // @[Mux.scala 46:19:@9604.4]
  wire [7:0] _T_10863; // @[Mux.scala 46:16:@9605.4]
  wire  _T_10864; // @[Mux.scala 46:19:@9606.4]
  wire [7:0] _T_10865; // @[Mux.scala 46:16:@9607.4]
  wire  _T_10866; // @[Mux.scala 46:19:@9608.4]
  wire [7:0] _T_10867; // @[Mux.scala 46:16:@9609.4]
  wire  _T_10868; // @[Mux.scala 46:19:@9610.4]
  wire [7:0] _T_10869; // @[Mux.scala 46:16:@9611.4]
  wire  _T_10870; // @[Mux.scala 46:19:@9612.4]
  wire [7:0] _T_10871; // @[Mux.scala 46:16:@9613.4]
  wire  _T_10872; // @[Mux.scala 46:19:@9614.4]
  wire [7:0] _T_10873; // @[Mux.scala 46:16:@9615.4]
  wire  _T_10874; // @[Mux.scala 46:19:@9616.4]
  wire [7:0] _T_10875; // @[Mux.scala 46:16:@9617.4]
  wire  _T_10876; // @[Mux.scala 46:19:@9618.4]
  wire [7:0] _T_10877; // @[Mux.scala 46:16:@9619.4]
  wire  _T_10878; // @[Mux.scala 46:19:@9620.4]
  wire [7:0] _T_10879; // @[Mux.scala 46:16:@9621.4]
  wire  _T_10880; // @[Mux.scala 46:19:@9622.4]
  wire [7:0] _T_10881; // @[Mux.scala 46:16:@9623.4]
  wire  _T_10882; // @[Mux.scala 46:19:@9624.4]
  wire [7:0] _T_10883; // @[Mux.scala 46:16:@9625.4]
  wire  _T_10884; // @[Mux.scala 46:19:@9626.4]
  wire [7:0] _T_10885; // @[Mux.scala 46:16:@9627.4]
  wire  _T_10905; // @[Mux.scala 46:19:@9629.4]
  wire [7:0] _T_10906; // @[Mux.scala 46:16:@9630.4]
  wire  _T_10907; // @[Mux.scala 46:19:@9631.4]
  wire [7:0] _T_10908; // @[Mux.scala 46:16:@9632.4]
  wire  _T_10909; // @[Mux.scala 46:19:@9633.4]
  wire [7:0] _T_10910; // @[Mux.scala 46:16:@9634.4]
  wire  _T_10911; // @[Mux.scala 46:19:@9635.4]
  wire [7:0] _T_10912; // @[Mux.scala 46:16:@9636.4]
  wire  _T_10913; // @[Mux.scala 46:19:@9637.4]
  wire [7:0] _T_10914; // @[Mux.scala 46:16:@9638.4]
  wire  _T_10915; // @[Mux.scala 46:19:@9639.4]
  wire [7:0] _T_10916; // @[Mux.scala 46:16:@9640.4]
  wire  _T_10917; // @[Mux.scala 46:19:@9641.4]
  wire [7:0] _T_10918; // @[Mux.scala 46:16:@9642.4]
  wire  _T_10919; // @[Mux.scala 46:19:@9643.4]
  wire [7:0] _T_10920; // @[Mux.scala 46:16:@9644.4]
  wire  _T_10921; // @[Mux.scala 46:19:@9645.4]
  wire [7:0] _T_10922; // @[Mux.scala 46:16:@9646.4]
  wire  _T_10923; // @[Mux.scala 46:19:@9647.4]
  wire [7:0] _T_10924; // @[Mux.scala 46:16:@9648.4]
  wire  _T_10925; // @[Mux.scala 46:19:@9649.4]
  wire [7:0] _T_10926; // @[Mux.scala 46:16:@9650.4]
  wire  _T_10927; // @[Mux.scala 46:19:@9651.4]
  wire [7:0] _T_10928; // @[Mux.scala 46:16:@9652.4]
  wire  _T_10929; // @[Mux.scala 46:19:@9653.4]
  wire [7:0] _T_10930; // @[Mux.scala 46:16:@9654.4]
  wire  _T_10931; // @[Mux.scala 46:19:@9655.4]
  wire [7:0] _T_10932; // @[Mux.scala 46:16:@9656.4]
  wire  _T_10933; // @[Mux.scala 46:19:@9657.4]
  wire [7:0] _T_10934; // @[Mux.scala 46:16:@9658.4]
  wire  _T_10935; // @[Mux.scala 46:19:@9659.4]
  wire [7:0] _T_10936; // @[Mux.scala 46:16:@9660.4]
  wire  _T_10937; // @[Mux.scala 46:19:@9661.4]
  wire [7:0] _T_10938; // @[Mux.scala 46:16:@9662.4]
  wire  _T_10939; // @[Mux.scala 46:19:@9663.4]
  wire [7:0] _T_10940; // @[Mux.scala 46:16:@9664.4]
  wire  _T_10961; // @[Mux.scala 46:19:@9666.4]
  wire [7:0] _T_10962; // @[Mux.scala 46:16:@9667.4]
  wire  _T_10963; // @[Mux.scala 46:19:@9668.4]
  wire [7:0] _T_10964; // @[Mux.scala 46:16:@9669.4]
  wire  _T_10965; // @[Mux.scala 46:19:@9670.4]
  wire [7:0] _T_10966; // @[Mux.scala 46:16:@9671.4]
  wire  _T_10967; // @[Mux.scala 46:19:@9672.4]
  wire [7:0] _T_10968; // @[Mux.scala 46:16:@9673.4]
  wire  _T_10969; // @[Mux.scala 46:19:@9674.4]
  wire [7:0] _T_10970; // @[Mux.scala 46:16:@9675.4]
  wire  _T_10971; // @[Mux.scala 46:19:@9676.4]
  wire [7:0] _T_10972; // @[Mux.scala 46:16:@9677.4]
  wire  _T_10973; // @[Mux.scala 46:19:@9678.4]
  wire [7:0] _T_10974; // @[Mux.scala 46:16:@9679.4]
  wire  _T_10975; // @[Mux.scala 46:19:@9680.4]
  wire [7:0] _T_10976; // @[Mux.scala 46:16:@9681.4]
  wire  _T_10977; // @[Mux.scala 46:19:@9682.4]
  wire [7:0] _T_10978; // @[Mux.scala 46:16:@9683.4]
  wire  _T_10979; // @[Mux.scala 46:19:@9684.4]
  wire [7:0] _T_10980; // @[Mux.scala 46:16:@9685.4]
  wire  _T_10981; // @[Mux.scala 46:19:@9686.4]
  wire [7:0] _T_10982; // @[Mux.scala 46:16:@9687.4]
  wire  _T_10983; // @[Mux.scala 46:19:@9688.4]
  wire [7:0] _T_10984; // @[Mux.scala 46:16:@9689.4]
  wire  _T_10985; // @[Mux.scala 46:19:@9690.4]
  wire [7:0] _T_10986; // @[Mux.scala 46:16:@9691.4]
  wire  _T_10987; // @[Mux.scala 46:19:@9692.4]
  wire [7:0] _T_10988; // @[Mux.scala 46:16:@9693.4]
  wire  _T_10989; // @[Mux.scala 46:19:@9694.4]
  wire [7:0] _T_10990; // @[Mux.scala 46:16:@9695.4]
  wire  _T_10991; // @[Mux.scala 46:19:@9696.4]
  wire [7:0] _T_10992; // @[Mux.scala 46:16:@9697.4]
  wire  _T_10993; // @[Mux.scala 46:19:@9698.4]
  wire [7:0] _T_10994; // @[Mux.scala 46:16:@9699.4]
  wire  _T_10995; // @[Mux.scala 46:19:@9700.4]
  wire [7:0] _T_10996; // @[Mux.scala 46:16:@9701.4]
  wire  _T_10997; // @[Mux.scala 46:19:@9702.4]
  wire [7:0] _T_10998; // @[Mux.scala 46:16:@9703.4]
  wire  _T_11020; // @[Mux.scala 46:19:@9705.4]
  wire [7:0] _T_11021; // @[Mux.scala 46:16:@9706.4]
  wire  _T_11022; // @[Mux.scala 46:19:@9707.4]
  wire [7:0] _T_11023; // @[Mux.scala 46:16:@9708.4]
  wire  _T_11024; // @[Mux.scala 46:19:@9709.4]
  wire [7:0] _T_11025; // @[Mux.scala 46:16:@9710.4]
  wire  _T_11026; // @[Mux.scala 46:19:@9711.4]
  wire [7:0] _T_11027; // @[Mux.scala 46:16:@9712.4]
  wire  _T_11028; // @[Mux.scala 46:19:@9713.4]
  wire [7:0] _T_11029; // @[Mux.scala 46:16:@9714.4]
  wire  _T_11030; // @[Mux.scala 46:19:@9715.4]
  wire [7:0] _T_11031; // @[Mux.scala 46:16:@9716.4]
  wire  _T_11032; // @[Mux.scala 46:19:@9717.4]
  wire [7:0] _T_11033; // @[Mux.scala 46:16:@9718.4]
  wire  _T_11034; // @[Mux.scala 46:19:@9719.4]
  wire [7:0] _T_11035; // @[Mux.scala 46:16:@9720.4]
  wire  _T_11036; // @[Mux.scala 46:19:@9721.4]
  wire [7:0] _T_11037; // @[Mux.scala 46:16:@9722.4]
  wire  _T_11038; // @[Mux.scala 46:19:@9723.4]
  wire [7:0] _T_11039; // @[Mux.scala 46:16:@9724.4]
  wire  _T_11040; // @[Mux.scala 46:19:@9725.4]
  wire [7:0] _T_11041; // @[Mux.scala 46:16:@9726.4]
  wire  _T_11042; // @[Mux.scala 46:19:@9727.4]
  wire [7:0] _T_11043; // @[Mux.scala 46:16:@9728.4]
  wire  _T_11044; // @[Mux.scala 46:19:@9729.4]
  wire [7:0] _T_11045; // @[Mux.scala 46:16:@9730.4]
  wire  _T_11046; // @[Mux.scala 46:19:@9731.4]
  wire [7:0] _T_11047; // @[Mux.scala 46:16:@9732.4]
  wire  _T_11048; // @[Mux.scala 46:19:@9733.4]
  wire [7:0] _T_11049; // @[Mux.scala 46:16:@9734.4]
  wire  _T_11050; // @[Mux.scala 46:19:@9735.4]
  wire [7:0] _T_11051; // @[Mux.scala 46:16:@9736.4]
  wire  _T_11052; // @[Mux.scala 46:19:@9737.4]
  wire [7:0] _T_11053; // @[Mux.scala 46:16:@9738.4]
  wire  _T_11054; // @[Mux.scala 46:19:@9739.4]
  wire [7:0] _T_11055; // @[Mux.scala 46:16:@9740.4]
  wire  _T_11056; // @[Mux.scala 46:19:@9741.4]
  wire [7:0] _T_11057; // @[Mux.scala 46:16:@9742.4]
  wire  _T_11058; // @[Mux.scala 46:19:@9743.4]
  wire [7:0] _T_11059; // @[Mux.scala 46:16:@9744.4]
  wire  _T_11082; // @[Mux.scala 46:19:@9746.4]
  wire [7:0] _T_11083; // @[Mux.scala 46:16:@9747.4]
  wire  _T_11084; // @[Mux.scala 46:19:@9748.4]
  wire [7:0] _T_11085; // @[Mux.scala 46:16:@9749.4]
  wire  _T_11086; // @[Mux.scala 46:19:@9750.4]
  wire [7:0] _T_11087; // @[Mux.scala 46:16:@9751.4]
  wire  _T_11088; // @[Mux.scala 46:19:@9752.4]
  wire [7:0] _T_11089; // @[Mux.scala 46:16:@9753.4]
  wire  _T_11090; // @[Mux.scala 46:19:@9754.4]
  wire [7:0] _T_11091; // @[Mux.scala 46:16:@9755.4]
  wire  _T_11092; // @[Mux.scala 46:19:@9756.4]
  wire [7:0] _T_11093; // @[Mux.scala 46:16:@9757.4]
  wire  _T_11094; // @[Mux.scala 46:19:@9758.4]
  wire [7:0] _T_11095; // @[Mux.scala 46:16:@9759.4]
  wire  _T_11096; // @[Mux.scala 46:19:@9760.4]
  wire [7:0] _T_11097; // @[Mux.scala 46:16:@9761.4]
  wire  _T_11098; // @[Mux.scala 46:19:@9762.4]
  wire [7:0] _T_11099; // @[Mux.scala 46:16:@9763.4]
  wire  _T_11100; // @[Mux.scala 46:19:@9764.4]
  wire [7:0] _T_11101; // @[Mux.scala 46:16:@9765.4]
  wire  _T_11102; // @[Mux.scala 46:19:@9766.4]
  wire [7:0] _T_11103; // @[Mux.scala 46:16:@9767.4]
  wire  _T_11104; // @[Mux.scala 46:19:@9768.4]
  wire [7:0] _T_11105; // @[Mux.scala 46:16:@9769.4]
  wire  _T_11106; // @[Mux.scala 46:19:@9770.4]
  wire [7:0] _T_11107; // @[Mux.scala 46:16:@9771.4]
  wire  _T_11108; // @[Mux.scala 46:19:@9772.4]
  wire [7:0] _T_11109; // @[Mux.scala 46:16:@9773.4]
  wire  _T_11110; // @[Mux.scala 46:19:@9774.4]
  wire [7:0] _T_11111; // @[Mux.scala 46:16:@9775.4]
  wire  _T_11112; // @[Mux.scala 46:19:@9776.4]
  wire [7:0] _T_11113; // @[Mux.scala 46:16:@9777.4]
  wire  _T_11114; // @[Mux.scala 46:19:@9778.4]
  wire [7:0] _T_11115; // @[Mux.scala 46:16:@9779.4]
  wire  _T_11116; // @[Mux.scala 46:19:@9780.4]
  wire [7:0] _T_11117; // @[Mux.scala 46:16:@9781.4]
  wire  _T_11118; // @[Mux.scala 46:19:@9782.4]
  wire [7:0] _T_11119; // @[Mux.scala 46:16:@9783.4]
  wire  _T_11120; // @[Mux.scala 46:19:@9784.4]
  wire [7:0] _T_11121; // @[Mux.scala 46:16:@9785.4]
  wire  _T_11122; // @[Mux.scala 46:19:@9786.4]
  wire [7:0] _T_11123; // @[Mux.scala 46:16:@9787.4]
  wire  _T_11147; // @[Mux.scala 46:19:@9789.4]
  wire [7:0] _T_11148; // @[Mux.scala 46:16:@9790.4]
  wire  _T_11149; // @[Mux.scala 46:19:@9791.4]
  wire [7:0] _T_11150; // @[Mux.scala 46:16:@9792.4]
  wire  _T_11151; // @[Mux.scala 46:19:@9793.4]
  wire [7:0] _T_11152; // @[Mux.scala 46:16:@9794.4]
  wire  _T_11153; // @[Mux.scala 46:19:@9795.4]
  wire [7:0] _T_11154; // @[Mux.scala 46:16:@9796.4]
  wire  _T_11155; // @[Mux.scala 46:19:@9797.4]
  wire [7:0] _T_11156; // @[Mux.scala 46:16:@9798.4]
  wire  _T_11157; // @[Mux.scala 46:19:@9799.4]
  wire [7:0] _T_11158; // @[Mux.scala 46:16:@9800.4]
  wire  _T_11159; // @[Mux.scala 46:19:@9801.4]
  wire [7:0] _T_11160; // @[Mux.scala 46:16:@9802.4]
  wire  _T_11161; // @[Mux.scala 46:19:@9803.4]
  wire [7:0] _T_11162; // @[Mux.scala 46:16:@9804.4]
  wire  _T_11163; // @[Mux.scala 46:19:@9805.4]
  wire [7:0] _T_11164; // @[Mux.scala 46:16:@9806.4]
  wire  _T_11165; // @[Mux.scala 46:19:@9807.4]
  wire [7:0] _T_11166; // @[Mux.scala 46:16:@9808.4]
  wire  _T_11167; // @[Mux.scala 46:19:@9809.4]
  wire [7:0] _T_11168; // @[Mux.scala 46:16:@9810.4]
  wire  _T_11169; // @[Mux.scala 46:19:@9811.4]
  wire [7:0] _T_11170; // @[Mux.scala 46:16:@9812.4]
  wire  _T_11171; // @[Mux.scala 46:19:@9813.4]
  wire [7:0] _T_11172; // @[Mux.scala 46:16:@9814.4]
  wire  _T_11173; // @[Mux.scala 46:19:@9815.4]
  wire [7:0] _T_11174; // @[Mux.scala 46:16:@9816.4]
  wire  _T_11175; // @[Mux.scala 46:19:@9817.4]
  wire [7:0] _T_11176; // @[Mux.scala 46:16:@9818.4]
  wire  _T_11177; // @[Mux.scala 46:19:@9819.4]
  wire [7:0] _T_11178; // @[Mux.scala 46:16:@9820.4]
  wire  _T_11179; // @[Mux.scala 46:19:@9821.4]
  wire [7:0] _T_11180; // @[Mux.scala 46:16:@9822.4]
  wire  _T_11181; // @[Mux.scala 46:19:@9823.4]
  wire [7:0] _T_11182; // @[Mux.scala 46:16:@9824.4]
  wire  _T_11183; // @[Mux.scala 46:19:@9825.4]
  wire [7:0] _T_11184; // @[Mux.scala 46:16:@9826.4]
  wire  _T_11185; // @[Mux.scala 46:19:@9827.4]
  wire [7:0] _T_11186; // @[Mux.scala 46:16:@9828.4]
  wire  _T_11187; // @[Mux.scala 46:19:@9829.4]
  wire [7:0] _T_11188; // @[Mux.scala 46:16:@9830.4]
  wire  _T_11189; // @[Mux.scala 46:19:@9831.4]
  wire [7:0] _T_11190; // @[Mux.scala 46:16:@9832.4]
  wire  _T_11215; // @[Mux.scala 46:19:@9834.4]
  wire [7:0] _T_11216; // @[Mux.scala 46:16:@9835.4]
  wire  _T_11217; // @[Mux.scala 46:19:@9836.4]
  wire [7:0] _T_11218; // @[Mux.scala 46:16:@9837.4]
  wire  _T_11219; // @[Mux.scala 46:19:@9838.4]
  wire [7:0] _T_11220; // @[Mux.scala 46:16:@9839.4]
  wire  _T_11221; // @[Mux.scala 46:19:@9840.4]
  wire [7:0] _T_11222; // @[Mux.scala 46:16:@9841.4]
  wire  _T_11223; // @[Mux.scala 46:19:@9842.4]
  wire [7:0] _T_11224; // @[Mux.scala 46:16:@9843.4]
  wire  _T_11225; // @[Mux.scala 46:19:@9844.4]
  wire [7:0] _T_11226; // @[Mux.scala 46:16:@9845.4]
  wire  _T_11227; // @[Mux.scala 46:19:@9846.4]
  wire [7:0] _T_11228; // @[Mux.scala 46:16:@9847.4]
  wire  _T_11229; // @[Mux.scala 46:19:@9848.4]
  wire [7:0] _T_11230; // @[Mux.scala 46:16:@9849.4]
  wire  _T_11231; // @[Mux.scala 46:19:@9850.4]
  wire [7:0] _T_11232; // @[Mux.scala 46:16:@9851.4]
  wire  _T_11233; // @[Mux.scala 46:19:@9852.4]
  wire [7:0] _T_11234; // @[Mux.scala 46:16:@9853.4]
  wire  _T_11235; // @[Mux.scala 46:19:@9854.4]
  wire [7:0] _T_11236; // @[Mux.scala 46:16:@9855.4]
  wire  _T_11237; // @[Mux.scala 46:19:@9856.4]
  wire [7:0] _T_11238; // @[Mux.scala 46:16:@9857.4]
  wire  _T_11239; // @[Mux.scala 46:19:@9858.4]
  wire [7:0] _T_11240; // @[Mux.scala 46:16:@9859.4]
  wire  _T_11241; // @[Mux.scala 46:19:@9860.4]
  wire [7:0] _T_11242; // @[Mux.scala 46:16:@9861.4]
  wire  _T_11243; // @[Mux.scala 46:19:@9862.4]
  wire [7:0] _T_11244; // @[Mux.scala 46:16:@9863.4]
  wire  _T_11245; // @[Mux.scala 46:19:@9864.4]
  wire [7:0] _T_11246; // @[Mux.scala 46:16:@9865.4]
  wire  _T_11247; // @[Mux.scala 46:19:@9866.4]
  wire [7:0] _T_11248; // @[Mux.scala 46:16:@9867.4]
  wire  _T_11249; // @[Mux.scala 46:19:@9868.4]
  wire [7:0] _T_11250; // @[Mux.scala 46:16:@9869.4]
  wire  _T_11251; // @[Mux.scala 46:19:@9870.4]
  wire [7:0] _T_11252; // @[Mux.scala 46:16:@9871.4]
  wire  _T_11253; // @[Mux.scala 46:19:@9872.4]
  wire [7:0] _T_11254; // @[Mux.scala 46:16:@9873.4]
  wire  _T_11255; // @[Mux.scala 46:19:@9874.4]
  wire [7:0] _T_11256; // @[Mux.scala 46:16:@9875.4]
  wire  _T_11257; // @[Mux.scala 46:19:@9876.4]
  wire [7:0] _T_11258; // @[Mux.scala 46:16:@9877.4]
  wire  _T_11259; // @[Mux.scala 46:19:@9878.4]
  wire [7:0] _T_11260; // @[Mux.scala 46:16:@9879.4]
  wire  _T_11286; // @[Mux.scala 46:19:@9881.4]
  wire [7:0] _T_11287; // @[Mux.scala 46:16:@9882.4]
  wire  _T_11288; // @[Mux.scala 46:19:@9883.4]
  wire [7:0] _T_11289; // @[Mux.scala 46:16:@9884.4]
  wire  _T_11290; // @[Mux.scala 46:19:@9885.4]
  wire [7:0] _T_11291; // @[Mux.scala 46:16:@9886.4]
  wire  _T_11292; // @[Mux.scala 46:19:@9887.4]
  wire [7:0] _T_11293; // @[Mux.scala 46:16:@9888.4]
  wire  _T_11294; // @[Mux.scala 46:19:@9889.4]
  wire [7:0] _T_11295; // @[Mux.scala 46:16:@9890.4]
  wire  _T_11296; // @[Mux.scala 46:19:@9891.4]
  wire [7:0] _T_11297; // @[Mux.scala 46:16:@9892.4]
  wire  _T_11298; // @[Mux.scala 46:19:@9893.4]
  wire [7:0] _T_11299; // @[Mux.scala 46:16:@9894.4]
  wire  _T_11300; // @[Mux.scala 46:19:@9895.4]
  wire [7:0] _T_11301; // @[Mux.scala 46:16:@9896.4]
  wire  _T_11302; // @[Mux.scala 46:19:@9897.4]
  wire [7:0] _T_11303; // @[Mux.scala 46:16:@9898.4]
  wire  _T_11304; // @[Mux.scala 46:19:@9899.4]
  wire [7:0] _T_11305; // @[Mux.scala 46:16:@9900.4]
  wire  _T_11306; // @[Mux.scala 46:19:@9901.4]
  wire [7:0] _T_11307; // @[Mux.scala 46:16:@9902.4]
  wire  _T_11308; // @[Mux.scala 46:19:@9903.4]
  wire [7:0] _T_11309; // @[Mux.scala 46:16:@9904.4]
  wire  _T_11310; // @[Mux.scala 46:19:@9905.4]
  wire [7:0] _T_11311; // @[Mux.scala 46:16:@9906.4]
  wire  _T_11312; // @[Mux.scala 46:19:@9907.4]
  wire [7:0] _T_11313; // @[Mux.scala 46:16:@9908.4]
  wire  _T_11314; // @[Mux.scala 46:19:@9909.4]
  wire [7:0] _T_11315; // @[Mux.scala 46:16:@9910.4]
  wire  _T_11316; // @[Mux.scala 46:19:@9911.4]
  wire [7:0] _T_11317; // @[Mux.scala 46:16:@9912.4]
  wire  _T_11318; // @[Mux.scala 46:19:@9913.4]
  wire [7:0] _T_11319; // @[Mux.scala 46:16:@9914.4]
  wire  _T_11320; // @[Mux.scala 46:19:@9915.4]
  wire [7:0] _T_11321; // @[Mux.scala 46:16:@9916.4]
  wire  _T_11322; // @[Mux.scala 46:19:@9917.4]
  wire [7:0] _T_11323; // @[Mux.scala 46:16:@9918.4]
  wire  _T_11324; // @[Mux.scala 46:19:@9919.4]
  wire [7:0] _T_11325; // @[Mux.scala 46:16:@9920.4]
  wire  _T_11326; // @[Mux.scala 46:19:@9921.4]
  wire [7:0] _T_11327; // @[Mux.scala 46:16:@9922.4]
  wire  _T_11328; // @[Mux.scala 46:19:@9923.4]
  wire [7:0] _T_11329; // @[Mux.scala 46:16:@9924.4]
  wire  _T_11330; // @[Mux.scala 46:19:@9925.4]
  wire [7:0] _T_11331; // @[Mux.scala 46:16:@9926.4]
  wire  _T_11332; // @[Mux.scala 46:19:@9927.4]
  wire [7:0] _T_11333; // @[Mux.scala 46:16:@9928.4]
  wire  _T_11360; // @[Mux.scala 46:19:@9930.4]
  wire [7:0] _T_11361; // @[Mux.scala 46:16:@9931.4]
  wire  _T_11362; // @[Mux.scala 46:19:@9932.4]
  wire [7:0] _T_11363; // @[Mux.scala 46:16:@9933.4]
  wire  _T_11364; // @[Mux.scala 46:19:@9934.4]
  wire [7:0] _T_11365; // @[Mux.scala 46:16:@9935.4]
  wire  _T_11366; // @[Mux.scala 46:19:@9936.4]
  wire [7:0] _T_11367; // @[Mux.scala 46:16:@9937.4]
  wire  _T_11368; // @[Mux.scala 46:19:@9938.4]
  wire [7:0] _T_11369; // @[Mux.scala 46:16:@9939.4]
  wire  _T_11370; // @[Mux.scala 46:19:@9940.4]
  wire [7:0] _T_11371; // @[Mux.scala 46:16:@9941.4]
  wire  _T_11372; // @[Mux.scala 46:19:@9942.4]
  wire [7:0] _T_11373; // @[Mux.scala 46:16:@9943.4]
  wire  _T_11374; // @[Mux.scala 46:19:@9944.4]
  wire [7:0] _T_11375; // @[Mux.scala 46:16:@9945.4]
  wire  _T_11376; // @[Mux.scala 46:19:@9946.4]
  wire [7:0] _T_11377; // @[Mux.scala 46:16:@9947.4]
  wire  _T_11378; // @[Mux.scala 46:19:@9948.4]
  wire [7:0] _T_11379; // @[Mux.scala 46:16:@9949.4]
  wire  _T_11380; // @[Mux.scala 46:19:@9950.4]
  wire [7:0] _T_11381; // @[Mux.scala 46:16:@9951.4]
  wire  _T_11382; // @[Mux.scala 46:19:@9952.4]
  wire [7:0] _T_11383; // @[Mux.scala 46:16:@9953.4]
  wire  _T_11384; // @[Mux.scala 46:19:@9954.4]
  wire [7:0] _T_11385; // @[Mux.scala 46:16:@9955.4]
  wire  _T_11386; // @[Mux.scala 46:19:@9956.4]
  wire [7:0] _T_11387; // @[Mux.scala 46:16:@9957.4]
  wire  _T_11388; // @[Mux.scala 46:19:@9958.4]
  wire [7:0] _T_11389; // @[Mux.scala 46:16:@9959.4]
  wire  _T_11390; // @[Mux.scala 46:19:@9960.4]
  wire [7:0] _T_11391; // @[Mux.scala 46:16:@9961.4]
  wire  _T_11392; // @[Mux.scala 46:19:@9962.4]
  wire [7:0] _T_11393; // @[Mux.scala 46:16:@9963.4]
  wire  _T_11394; // @[Mux.scala 46:19:@9964.4]
  wire [7:0] _T_11395; // @[Mux.scala 46:16:@9965.4]
  wire  _T_11396; // @[Mux.scala 46:19:@9966.4]
  wire [7:0] _T_11397; // @[Mux.scala 46:16:@9967.4]
  wire  _T_11398; // @[Mux.scala 46:19:@9968.4]
  wire [7:0] _T_11399; // @[Mux.scala 46:16:@9969.4]
  wire  _T_11400; // @[Mux.scala 46:19:@9970.4]
  wire [7:0] _T_11401; // @[Mux.scala 46:16:@9971.4]
  wire  _T_11402; // @[Mux.scala 46:19:@9972.4]
  wire [7:0] _T_11403; // @[Mux.scala 46:16:@9973.4]
  wire  _T_11404; // @[Mux.scala 46:19:@9974.4]
  wire [7:0] _T_11405; // @[Mux.scala 46:16:@9975.4]
  wire  _T_11406; // @[Mux.scala 46:19:@9976.4]
  wire [7:0] _T_11407; // @[Mux.scala 46:16:@9977.4]
  wire  _T_11408; // @[Mux.scala 46:19:@9978.4]
  wire [7:0] _T_11409; // @[Mux.scala 46:16:@9979.4]
  wire  _T_11437; // @[Mux.scala 46:19:@9981.4]
  wire [7:0] _T_11438; // @[Mux.scala 46:16:@9982.4]
  wire  _T_11439; // @[Mux.scala 46:19:@9983.4]
  wire [7:0] _T_11440; // @[Mux.scala 46:16:@9984.4]
  wire  _T_11441; // @[Mux.scala 46:19:@9985.4]
  wire [7:0] _T_11442; // @[Mux.scala 46:16:@9986.4]
  wire  _T_11443; // @[Mux.scala 46:19:@9987.4]
  wire [7:0] _T_11444; // @[Mux.scala 46:16:@9988.4]
  wire  _T_11445; // @[Mux.scala 46:19:@9989.4]
  wire [7:0] _T_11446; // @[Mux.scala 46:16:@9990.4]
  wire  _T_11447; // @[Mux.scala 46:19:@9991.4]
  wire [7:0] _T_11448; // @[Mux.scala 46:16:@9992.4]
  wire  _T_11449; // @[Mux.scala 46:19:@9993.4]
  wire [7:0] _T_11450; // @[Mux.scala 46:16:@9994.4]
  wire  _T_11451; // @[Mux.scala 46:19:@9995.4]
  wire [7:0] _T_11452; // @[Mux.scala 46:16:@9996.4]
  wire  _T_11453; // @[Mux.scala 46:19:@9997.4]
  wire [7:0] _T_11454; // @[Mux.scala 46:16:@9998.4]
  wire  _T_11455; // @[Mux.scala 46:19:@9999.4]
  wire [7:0] _T_11456; // @[Mux.scala 46:16:@10000.4]
  wire  _T_11457; // @[Mux.scala 46:19:@10001.4]
  wire [7:0] _T_11458; // @[Mux.scala 46:16:@10002.4]
  wire  _T_11459; // @[Mux.scala 46:19:@10003.4]
  wire [7:0] _T_11460; // @[Mux.scala 46:16:@10004.4]
  wire  _T_11461; // @[Mux.scala 46:19:@10005.4]
  wire [7:0] _T_11462; // @[Mux.scala 46:16:@10006.4]
  wire  _T_11463; // @[Mux.scala 46:19:@10007.4]
  wire [7:0] _T_11464; // @[Mux.scala 46:16:@10008.4]
  wire  _T_11465; // @[Mux.scala 46:19:@10009.4]
  wire [7:0] _T_11466; // @[Mux.scala 46:16:@10010.4]
  wire  _T_11467; // @[Mux.scala 46:19:@10011.4]
  wire [7:0] _T_11468; // @[Mux.scala 46:16:@10012.4]
  wire  _T_11469; // @[Mux.scala 46:19:@10013.4]
  wire [7:0] _T_11470; // @[Mux.scala 46:16:@10014.4]
  wire  _T_11471; // @[Mux.scala 46:19:@10015.4]
  wire [7:0] _T_11472; // @[Mux.scala 46:16:@10016.4]
  wire  _T_11473; // @[Mux.scala 46:19:@10017.4]
  wire [7:0] _T_11474; // @[Mux.scala 46:16:@10018.4]
  wire  _T_11475; // @[Mux.scala 46:19:@10019.4]
  wire [7:0] _T_11476; // @[Mux.scala 46:16:@10020.4]
  wire  _T_11477; // @[Mux.scala 46:19:@10021.4]
  wire [7:0] _T_11478; // @[Mux.scala 46:16:@10022.4]
  wire  _T_11479; // @[Mux.scala 46:19:@10023.4]
  wire [7:0] _T_11480; // @[Mux.scala 46:16:@10024.4]
  wire  _T_11481; // @[Mux.scala 46:19:@10025.4]
  wire [7:0] _T_11482; // @[Mux.scala 46:16:@10026.4]
  wire  _T_11483; // @[Mux.scala 46:19:@10027.4]
  wire [7:0] _T_11484; // @[Mux.scala 46:16:@10028.4]
  wire  _T_11485; // @[Mux.scala 46:19:@10029.4]
  wire [7:0] _T_11486; // @[Mux.scala 46:16:@10030.4]
  wire  _T_11487; // @[Mux.scala 46:19:@10031.4]
  wire [7:0] _T_11488; // @[Mux.scala 46:16:@10032.4]
  wire  _T_11517; // @[Mux.scala 46:19:@10034.4]
  wire [7:0] _T_11518; // @[Mux.scala 46:16:@10035.4]
  wire  _T_11519; // @[Mux.scala 46:19:@10036.4]
  wire [7:0] _T_11520; // @[Mux.scala 46:16:@10037.4]
  wire  _T_11521; // @[Mux.scala 46:19:@10038.4]
  wire [7:0] _T_11522; // @[Mux.scala 46:16:@10039.4]
  wire  _T_11523; // @[Mux.scala 46:19:@10040.4]
  wire [7:0] _T_11524; // @[Mux.scala 46:16:@10041.4]
  wire  _T_11525; // @[Mux.scala 46:19:@10042.4]
  wire [7:0] _T_11526; // @[Mux.scala 46:16:@10043.4]
  wire  _T_11527; // @[Mux.scala 46:19:@10044.4]
  wire [7:0] _T_11528; // @[Mux.scala 46:16:@10045.4]
  wire  _T_11529; // @[Mux.scala 46:19:@10046.4]
  wire [7:0] _T_11530; // @[Mux.scala 46:16:@10047.4]
  wire  _T_11531; // @[Mux.scala 46:19:@10048.4]
  wire [7:0] _T_11532; // @[Mux.scala 46:16:@10049.4]
  wire  _T_11533; // @[Mux.scala 46:19:@10050.4]
  wire [7:0] _T_11534; // @[Mux.scala 46:16:@10051.4]
  wire  _T_11535; // @[Mux.scala 46:19:@10052.4]
  wire [7:0] _T_11536; // @[Mux.scala 46:16:@10053.4]
  wire  _T_11537; // @[Mux.scala 46:19:@10054.4]
  wire [7:0] _T_11538; // @[Mux.scala 46:16:@10055.4]
  wire  _T_11539; // @[Mux.scala 46:19:@10056.4]
  wire [7:0] _T_11540; // @[Mux.scala 46:16:@10057.4]
  wire  _T_11541; // @[Mux.scala 46:19:@10058.4]
  wire [7:0] _T_11542; // @[Mux.scala 46:16:@10059.4]
  wire  _T_11543; // @[Mux.scala 46:19:@10060.4]
  wire [7:0] _T_11544; // @[Mux.scala 46:16:@10061.4]
  wire  _T_11545; // @[Mux.scala 46:19:@10062.4]
  wire [7:0] _T_11546; // @[Mux.scala 46:16:@10063.4]
  wire  _T_11547; // @[Mux.scala 46:19:@10064.4]
  wire [7:0] _T_11548; // @[Mux.scala 46:16:@10065.4]
  wire  _T_11549; // @[Mux.scala 46:19:@10066.4]
  wire [7:0] _T_11550; // @[Mux.scala 46:16:@10067.4]
  wire  _T_11551; // @[Mux.scala 46:19:@10068.4]
  wire [7:0] _T_11552; // @[Mux.scala 46:16:@10069.4]
  wire  _T_11553; // @[Mux.scala 46:19:@10070.4]
  wire [7:0] _T_11554; // @[Mux.scala 46:16:@10071.4]
  wire  _T_11555; // @[Mux.scala 46:19:@10072.4]
  wire [7:0] _T_11556; // @[Mux.scala 46:16:@10073.4]
  wire  _T_11557; // @[Mux.scala 46:19:@10074.4]
  wire [7:0] _T_11558; // @[Mux.scala 46:16:@10075.4]
  wire  _T_11559; // @[Mux.scala 46:19:@10076.4]
  wire [7:0] _T_11560; // @[Mux.scala 46:16:@10077.4]
  wire  _T_11561; // @[Mux.scala 46:19:@10078.4]
  wire [7:0] _T_11562; // @[Mux.scala 46:16:@10079.4]
  wire  _T_11563; // @[Mux.scala 46:19:@10080.4]
  wire [7:0] _T_11564; // @[Mux.scala 46:16:@10081.4]
  wire  _T_11565; // @[Mux.scala 46:19:@10082.4]
  wire [7:0] _T_11566; // @[Mux.scala 46:16:@10083.4]
  wire  _T_11567; // @[Mux.scala 46:19:@10084.4]
  wire [7:0] _T_11568; // @[Mux.scala 46:16:@10085.4]
  wire  _T_11569; // @[Mux.scala 46:19:@10086.4]
  wire [7:0] _T_11570; // @[Mux.scala 46:16:@10087.4]
  wire  _T_11600; // @[Mux.scala 46:19:@10089.4]
  wire [7:0] _T_11601; // @[Mux.scala 46:16:@10090.4]
  wire  _T_11602; // @[Mux.scala 46:19:@10091.4]
  wire [7:0] _T_11603; // @[Mux.scala 46:16:@10092.4]
  wire  _T_11604; // @[Mux.scala 46:19:@10093.4]
  wire [7:0] _T_11605; // @[Mux.scala 46:16:@10094.4]
  wire  _T_11606; // @[Mux.scala 46:19:@10095.4]
  wire [7:0] _T_11607; // @[Mux.scala 46:16:@10096.4]
  wire  _T_11608; // @[Mux.scala 46:19:@10097.4]
  wire [7:0] _T_11609; // @[Mux.scala 46:16:@10098.4]
  wire  _T_11610; // @[Mux.scala 46:19:@10099.4]
  wire [7:0] _T_11611; // @[Mux.scala 46:16:@10100.4]
  wire  _T_11612; // @[Mux.scala 46:19:@10101.4]
  wire [7:0] _T_11613; // @[Mux.scala 46:16:@10102.4]
  wire  _T_11614; // @[Mux.scala 46:19:@10103.4]
  wire [7:0] _T_11615; // @[Mux.scala 46:16:@10104.4]
  wire  _T_11616; // @[Mux.scala 46:19:@10105.4]
  wire [7:0] _T_11617; // @[Mux.scala 46:16:@10106.4]
  wire  _T_11618; // @[Mux.scala 46:19:@10107.4]
  wire [7:0] _T_11619; // @[Mux.scala 46:16:@10108.4]
  wire  _T_11620; // @[Mux.scala 46:19:@10109.4]
  wire [7:0] _T_11621; // @[Mux.scala 46:16:@10110.4]
  wire  _T_11622; // @[Mux.scala 46:19:@10111.4]
  wire [7:0] _T_11623; // @[Mux.scala 46:16:@10112.4]
  wire  _T_11624; // @[Mux.scala 46:19:@10113.4]
  wire [7:0] _T_11625; // @[Mux.scala 46:16:@10114.4]
  wire  _T_11626; // @[Mux.scala 46:19:@10115.4]
  wire [7:0] _T_11627; // @[Mux.scala 46:16:@10116.4]
  wire  _T_11628; // @[Mux.scala 46:19:@10117.4]
  wire [7:0] _T_11629; // @[Mux.scala 46:16:@10118.4]
  wire  _T_11630; // @[Mux.scala 46:19:@10119.4]
  wire [7:0] _T_11631; // @[Mux.scala 46:16:@10120.4]
  wire  _T_11632; // @[Mux.scala 46:19:@10121.4]
  wire [7:0] _T_11633; // @[Mux.scala 46:16:@10122.4]
  wire  _T_11634; // @[Mux.scala 46:19:@10123.4]
  wire [7:0] _T_11635; // @[Mux.scala 46:16:@10124.4]
  wire  _T_11636; // @[Mux.scala 46:19:@10125.4]
  wire [7:0] _T_11637; // @[Mux.scala 46:16:@10126.4]
  wire  _T_11638; // @[Mux.scala 46:19:@10127.4]
  wire [7:0] _T_11639; // @[Mux.scala 46:16:@10128.4]
  wire  _T_11640; // @[Mux.scala 46:19:@10129.4]
  wire [7:0] _T_11641; // @[Mux.scala 46:16:@10130.4]
  wire  _T_11642; // @[Mux.scala 46:19:@10131.4]
  wire [7:0] _T_11643; // @[Mux.scala 46:16:@10132.4]
  wire  _T_11644; // @[Mux.scala 46:19:@10133.4]
  wire [7:0] _T_11645; // @[Mux.scala 46:16:@10134.4]
  wire  _T_11646; // @[Mux.scala 46:19:@10135.4]
  wire [7:0] _T_11647; // @[Mux.scala 46:16:@10136.4]
  wire  _T_11648; // @[Mux.scala 46:19:@10137.4]
  wire [7:0] _T_11649; // @[Mux.scala 46:16:@10138.4]
  wire  _T_11650; // @[Mux.scala 46:19:@10139.4]
  wire [7:0] _T_11651; // @[Mux.scala 46:16:@10140.4]
  wire  _T_11652; // @[Mux.scala 46:19:@10141.4]
  wire [7:0] _T_11653; // @[Mux.scala 46:16:@10142.4]
  wire  _T_11654; // @[Mux.scala 46:19:@10143.4]
  wire [7:0] _T_11655; // @[Mux.scala 46:16:@10144.4]
  wire  _T_11686; // @[Mux.scala 46:19:@10146.4]
  wire [7:0] _T_11687; // @[Mux.scala 46:16:@10147.4]
  wire  _T_11688; // @[Mux.scala 46:19:@10148.4]
  wire [7:0] _T_11689; // @[Mux.scala 46:16:@10149.4]
  wire  _T_11690; // @[Mux.scala 46:19:@10150.4]
  wire [7:0] _T_11691; // @[Mux.scala 46:16:@10151.4]
  wire  _T_11692; // @[Mux.scala 46:19:@10152.4]
  wire [7:0] _T_11693; // @[Mux.scala 46:16:@10153.4]
  wire  _T_11694; // @[Mux.scala 46:19:@10154.4]
  wire [7:0] _T_11695; // @[Mux.scala 46:16:@10155.4]
  wire  _T_11696; // @[Mux.scala 46:19:@10156.4]
  wire [7:0] _T_11697; // @[Mux.scala 46:16:@10157.4]
  wire  _T_11698; // @[Mux.scala 46:19:@10158.4]
  wire [7:0] _T_11699; // @[Mux.scala 46:16:@10159.4]
  wire  _T_11700; // @[Mux.scala 46:19:@10160.4]
  wire [7:0] _T_11701; // @[Mux.scala 46:16:@10161.4]
  wire  _T_11702; // @[Mux.scala 46:19:@10162.4]
  wire [7:0] _T_11703; // @[Mux.scala 46:16:@10163.4]
  wire  _T_11704; // @[Mux.scala 46:19:@10164.4]
  wire [7:0] _T_11705; // @[Mux.scala 46:16:@10165.4]
  wire  _T_11706; // @[Mux.scala 46:19:@10166.4]
  wire [7:0] _T_11707; // @[Mux.scala 46:16:@10167.4]
  wire  _T_11708; // @[Mux.scala 46:19:@10168.4]
  wire [7:0] _T_11709; // @[Mux.scala 46:16:@10169.4]
  wire  _T_11710; // @[Mux.scala 46:19:@10170.4]
  wire [7:0] _T_11711; // @[Mux.scala 46:16:@10171.4]
  wire  _T_11712; // @[Mux.scala 46:19:@10172.4]
  wire [7:0] _T_11713; // @[Mux.scala 46:16:@10173.4]
  wire  _T_11714; // @[Mux.scala 46:19:@10174.4]
  wire [7:0] _T_11715; // @[Mux.scala 46:16:@10175.4]
  wire  _T_11716; // @[Mux.scala 46:19:@10176.4]
  wire [7:0] _T_11717; // @[Mux.scala 46:16:@10177.4]
  wire  _T_11718; // @[Mux.scala 46:19:@10178.4]
  wire [7:0] _T_11719; // @[Mux.scala 46:16:@10179.4]
  wire  _T_11720; // @[Mux.scala 46:19:@10180.4]
  wire [7:0] _T_11721; // @[Mux.scala 46:16:@10181.4]
  wire  _T_11722; // @[Mux.scala 46:19:@10182.4]
  wire [7:0] _T_11723; // @[Mux.scala 46:16:@10183.4]
  wire  _T_11724; // @[Mux.scala 46:19:@10184.4]
  wire [7:0] _T_11725; // @[Mux.scala 46:16:@10185.4]
  wire  _T_11726; // @[Mux.scala 46:19:@10186.4]
  wire [7:0] _T_11727; // @[Mux.scala 46:16:@10187.4]
  wire  _T_11728; // @[Mux.scala 46:19:@10188.4]
  wire [7:0] _T_11729; // @[Mux.scala 46:16:@10189.4]
  wire  _T_11730; // @[Mux.scala 46:19:@10190.4]
  wire [7:0] _T_11731; // @[Mux.scala 46:16:@10191.4]
  wire  _T_11732; // @[Mux.scala 46:19:@10192.4]
  wire [7:0] _T_11733; // @[Mux.scala 46:16:@10193.4]
  wire  _T_11734; // @[Mux.scala 46:19:@10194.4]
  wire [7:0] _T_11735; // @[Mux.scala 46:16:@10195.4]
  wire  _T_11736; // @[Mux.scala 46:19:@10196.4]
  wire [7:0] _T_11737; // @[Mux.scala 46:16:@10197.4]
  wire  _T_11738; // @[Mux.scala 46:19:@10198.4]
  wire [7:0] _T_11739; // @[Mux.scala 46:16:@10199.4]
  wire  _T_11740; // @[Mux.scala 46:19:@10200.4]
  wire [7:0] _T_11741; // @[Mux.scala 46:16:@10201.4]
  wire  _T_11742; // @[Mux.scala 46:19:@10202.4]
  wire [7:0] _T_11743; // @[Mux.scala 46:16:@10203.4]
  wire  _T_11775; // @[Mux.scala 46:19:@10205.4]
  wire [7:0] _T_11776; // @[Mux.scala 46:16:@10206.4]
  wire  _T_11777; // @[Mux.scala 46:19:@10207.4]
  wire [7:0] _T_11778; // @[Mux.scala 46:16:@10208.4]
  wire  _T_11779; // @[Mux.scala 46:19:@10209.4]
  wire [7:0] _T_11780; // @[Mux.scala 46:16:@10210.4]
  wire  _T_11781; // @[Mux.scala 46:19:@10211.4]
  wire [7:0] _T_11782; // @[Mux.scala 46:16:@10212.4]
  wire  _T_11783; // @[Mux.scala 46:19:@10213.4]
  wire [7:0] _T_11784; // @[Mux.scala 46:16:@10214.4]
  wire  _T_11785; // @[Mux.scala 46:19:@10215.4]
  wire [7:0] _T_11786; // @[Mux.scala 46:16:@10216.4]
  wire  _T_11787; // @[Mux.scala 46:19:@10217.4]
  wire [7:0] _T_11788; // @[Mux.scala 46:16:@10218.4]
  wire  _T_11789; // @[Mux.scala 46:19:@10219.4]
  wire [7:0] _T_11790; // @[Mux.scala 46:16:@10220.4]
  wire  _T_11791; // @[Mux.scala 46:19:@10221.4]
  wire [7:0] _T_11792; // @[Mux.scala 46:16:@10222.4]
  wire  _T_11793; // @[Mux.scala 46:19:@10223.4]
  wire [7:0] _T_11794; // @[Mux.scala 46:16:@10224.4]
  wire  _T_11795; // @[Mux.scala 46:19:@10225.4]
  wire [7:0] _T_11796; // @[Mux.scala 46:16:@10226.4]
  wire  _T_11797; // @[Mux.scala 46:19:@10227.4]
  wire [7:0] _T_11798; // @[Mux.scala 46:16:@10228.4]
  wire  _T_11799; // @[Mux.scala 46:19:@10229.4]
  wire [7:0] _T_11800; // @[Mux.scala 46:16:@10230.4]
  wire  _T_11801; // @[Mux.scala 46:19:@10231.4]
  wire [7:0] _T_11802; // @[Mux.scala 46:16:@10232.4]
  wire  _T_11803; // @[Mux.scala 46:19:@10233.4]
  wire [7:0] _T_11804; // @[Mux.scala 46:16:@10234.4]
  wire  _T_11805; // @[Mux.scala 46:19:@10235.4]
  wire [7:0] _T_11806; // @[Mux.scala 46:16:@10236.4]
  wire  _T_11807; // @[Mux.scala 46:19:@10237.4]
  wire [7:0] _T_11808; // @[Mux.scala 46:16:@10238.4]
  wire  _T_11809; // @[Mux.scala 46:19:@10239.4]
  wire [7:0] _T_11810; // @[Mux.scala 46:16:@10240.4]
  wire  _T_11811; // @[Mux.scala 46:19:@10241.4]
  wire [7:0] _T_11812; // @[Mux.scala 46:16:@10242.4]
  wire  _T_11813; // @[Mux.scala 46:19:@10243.4]
  wire [7:0] _T_11814; // @[Mux.scala 46:16:@10244.4]
  wire  _T_11815; // @[Mux.scala 46:19:@10245.4]
  wire [7:0] _T_11816; // @[Mux.scala 46:16:@10246.4]
  wire  _T_11817; // @[Mux.scala 46:19:@10247.4]
  wire [7:0] _T_11818; // @[Mux.scala 46:16:@10248.4]
  wire  _T_11819; // @[Mux.scala 46:19:@10249.4]
  wire [7:0] _T_11820; // @[Mux.scala 46:16:@10250.4]
  wire  _T_11821; // @[Mux.scala 46:19:@10251.4]
  wire [7:0] _T_11822; // @[Mux.scala 46:16:@10252.4]
  wire  _T_11823; // @[Mux.scala 46:19:@10253.4]
  wire [7:0] _T_11824; // @[Mux.scala 46:16:@10254.4]
  wire  _T_11825; // @[Mux.scala 46:19:@10255.4]
  wire [7:0] _T_11826; // @[Mux.scala 46:16:@10256.4]
  wire  _T_11827; // @[Mux.scala 46:19:@10257.4]
  wire [7:0] _T_11828; // @[Mux.scala 46:16:@10258.4]
  wire  _T_11829; // @[Mux.scala 46:19:@10259.4]
  wire [7:0] _T_11830; // @[Mux.scala 46:16:@10260.4]
  wire  _T_11831; // @[Mux.scala 46:19:@10261.4]
  wire [7:0] _T_11832; // @[Mux.scala 46:16:@10262.4]
  wire  _T_11833; // @[Mux.scala 46:19:@10263.4]
  wire [7:0] _T_11834; // @[Mux.scala 46:16:@10264.4]
  wire  _T_11867; // @[Mux.scala 46:19:@10266.4]
  wire [7:0] _T_11868; // @[Mux.scala 46:16:@10267.4]
  wire  _T_11869; // @[Mux.scala 46:19:@10268.4]
  wire [7:0] _T_11870; // @[Mux.scala 46:16:@10269.4]
  wire  _T_11871; // @[Mux.scala 46:19:@10270.4]
  wire [7:0] _T_11872; // @[Mux.scala 46:16:@10271.4]
  wire  _T_11873; // @[Mux.scala 46:19:@10272.4]
  wire [7:0] _T_11874; // @[Mux.scala 46:16:@10273.4]
  wire  _T_11875; // @[Mux.scala 46:19:@10274.4]
  wire [7:0] _T_11876; // @[Mux.scala 46:16:@10275.4]
  wire  _T_11877; // @[Mux.scala 46:19:@10276.4]
  wire [7:0] _T_11878; // @[Mux.scala 46:16:@10277.4]
  wire  _T_11879; // @[Mux.scala 46:19:@10278.4]
  wire [7:0] _T_11880; // @[Mux.scala 46:16:@10279.4]
  wire  _T_11881; // @[Mux.scala 46:19:@10280.4]
  wire [7:0] _T_11882; // @[Mux.scala 46:16:@10281.4]
  wire  _T_11883; // @[Mux.scala 46:19:@10282.4]
  wire [7:0] _T_11884; // @[Mux.scala 46:16:@10283.4]
  wire  _T_11885; // @[Mux.scala 46:19:@10284.4]
  wire [7:0] _T_11886; // @[Mux.scala 46:16:@10285.4]
  wire  _T_11887; // @[Mux.scala 46:19:@10286.4]
  wire [7:0] _T_11888; // @[Mux.scala 46:16:@10287.4]
  wire  _T_11889; // @[Mux.scala 46:19:@10288.4]
  wire [7:0] _T_11890; // @[Mux.scala 46:16:@10289.4]
  wire  _T_11891; // @[Mux.scala 46:19:@10290.4]
  wire [7:0] _T_11892; // @[Mux.scala 46:16:@10291.4]
  wire  _T_11893; // @[Mux.scala 46:19:@10292.4]
  wire [7:0] _T_11894; // @[Mux.scala 46:16:@10293.4]
  wire  _T_11895; // @[Mux.scala 46:19:@10294.4]
  wire [7:0] _T_11896; // @[Mux.scala 46:16:@10295.4]
  wire  _T_11897; // @[Mux.scala 46:19:@10296.4]
  wire [7:0] _T_11898; // @[Mux.scala 46:16:@10297.4]
  wire  _T_11899; // @[Mux.scala 46:19:@10298.4]
  wire [7:0] _T_11900; // @[Mux.scala 46:16:@10299.4]
  wire  _T_11901; // @[Mux.scala 46:19:@10300.4]
  wire [7:0] _T_11902; // @[Mux.scala 46:16:@10301.4]
  wire  _T_11903; // @[Mux.scala 46:19:@10302.4]
  wire [7:0] _T_11904; // @[Mux.scala 46:16:@10303.4]
  wire  _T_11905; // @[Mux.scala 46:19:@10304.4]
  wire [7:0] _T_11906; // @[Mux.scala 46:16:@10305.4]
  wire  _T_11907; // @[Mux.scala 46:19:@10306.4]
  wire [7:0] _T_11908; // @[Mux.scala 46:16:@10307.4]
  wire  _T_11909; // @[Mux.scala 46:19:@10308.4]
  wire [7:0] _T_11910; // @[Mux.scala 46:16:@10309.4]
  wire  _T_11911; // @[Mux.scala 46:19:@10310.4]
  wire [7:0] _T_11912; // @[Mux.scala 46:16:@10311.4]
  wire  _T_11913; // @[Mux.scala 46:19:@10312.4]
  wire [7:0] _T_11914; // @[Mux.scala 46:16:@10313.4]
  wire  _T_11915; // @[Mux.scala 46:19:@10314.4]
  wire [7:0] _T_11916; // @[Mux.scala 46:16:@10315.4]
  wire  _T_11917; // @[Mux.scala 46:19:@10316.4]
  wire [7:0] _T_11918; // @[Mux.scala 46:16:@10317.4]
  wire  _T_11919; // @[Mux.scala 46:19:@10318.4]
  wire [7:0] _T_11920; // @[Mux.scala 46:16:@10319.4]
  wire  _T_11921; // @[Mux.scala 46:19:@10320.4]
  wire [7:0] _T_11922; // @[Mux.scala 46:16:@10321.4]
  wire  _T_11923; // @[Mux.scala 46:19:@10322.4]
  wire [7:0] _T_11924; // @[Mux.scala 46:16:@10323.4]
  wire  _T_11925; // @[Mux.scala 46:19:@10324.4]
  wire [7:0] _T_11926; // @[Mux.scala 46:16:@10325.4]
  wire  _T_11927; // @[Mux.scala 46:19:@10326.4]
  wire [7:0] _T_11928; // @[Mux.scala 46:16:@10327.4]
  wire  _T_11962; // @[Mux.scala 46:19:@10329.4]
  wire [7:0] _T_11963; // @[Mux.scala 46:16:@10330.4]
  wire  _T_11964; // @[Mux.scala 46:19:@10331.4]
  wire [7:0] _T_11965; // @[Mux.scala 46:16:@10332.4]
  wire  _T_11966; // @[Mux.scala 46:19:@10333.4]
  wire [7:0] _T_11967; // @[Mux.scala 46:16:@10334.4]
  wire  _T_11968; // @[Mux.scala 46:19:@10335.4]
  wire [7:0] _T_11969; // @[Mux.scala 46:16:@10336.4]
  wire  _T_11970; // @[Mux.scala 46:19:@10337.4]
  wire [7:0] _T_11971; // @[Mux.scala 46:16:@10338.4]
  wire  _T_11972; // @[Mux.scala 46:19:@10339.4]
  wire [7:0] _T_11973; // @[Mux.scala 46:16:@10340.4]
  wire  _T_11974; // @[Mux.scala 46:19:@10341.4]
  wire [7:0] _T_11975; // @[Mux.scala 46:16:@10342.4]
  wire  _T_11976; // @[Mux.scala 46:19:@10343.4]
  wire [7:0] _T_11977; // @[Mux.scala 46:16:@10344.4]
  wire  _T_11978; // @[Mux.scala 46:19:@10345.4]
  wire [7:0] _T_11979; // @[Mux.scala 46:16:@10346.4]
  wire  _T_11980; // @[Mux.scala 46:19:@10347.4]
  wire [7:0] _T_11981; // @[Mux.scala 46:16:@10348.4]
  wire  _T_11982; // @[Mux.scala 46:19:@10349.4]
  wire [7:0] _T_11983; // @[Mux.scala 46:16:@10350.4]
  wire  _T_11984; // @[Mux.scala 46:19:@10351.4]
  wire [7:0] _T_11985; // @[Mux.scala 46:16:@10352.4]
  wire  _T_11986; // @[Mux.scala 46:19:@10353.4]
  wire [7:0] _T_11987; // @[Mux.scala 46:16:@10354.4]
  wire  _T_11988; // @[Mux.scala 46:19:@10355.4]
  wire [7:0] _T_11989; // @[Mux.scala 46:16:@10356.4]
  wire  _T_11990; // @[Mux.scala 46:19:@10357.4]
  wire [7:0] _T_11991; // @[Mux.scala 46:16:@10358.4]
  wire  _T_11992; // @[Mux.scala 46:19:@10359.4]
  wire [7:0] _T_11993; // @[Mux.scala 46:16:@10360.4]
  wire  _T_11994; // @[Mux.scala 46:19:@10361.4]
  wire [7:0] _T_11995; // @[Mux.scala 46:16:@10362.4]
  wire  _T_11996; // @[Mux.scala 46:19:@10363.4]
  wire [7:0] _T_11997; // @[Mux.scala 46:16:@10364.4]
  wire  _T_11998; // @[Mux.scala 46:19:@10365.4]
  wire [7:0] _T_11999; // @[Mux.scala 46:16:@10366.4]
  wire  _T_12000; // @[Mux.scala 46:19:@10367.4]
  wire [7:0] _T_12001; // @[Mux.scala 46:16:@10368.4]
  wire  _T_12002; // @[Mux.scala 46:19:@10369.4]
  wire [7:0] _T_12003; // @[Mux.scala 46:16:@10370.4]
  wire  _T_12004; // @[Mux.scala 46:19:@10371.4]
  wire [7:0] _T_12005; // @[Mux.scala 46:16:@10372.4]
  wire  _T_12006; // @[Mux.scala 46:19:@10373.4]
  wire [7:0] _T_12007; // @[Mux.scala 46:16:@10374.4]
  wire  _T_12008; // @[Mux.scala 46:19:@10375.4]
  wire [7:0] _T_12009; // @[Mux.scala 46:16:@10376.4]
  wire  _T_12010; // @[Mux.scala 46:19:@10377.4]
  wire [7:0] _T_12011; // @[Mux.scala 46:16:@10378.4]
  wire  _T_12012; // @[Mux.scala 46:19:@10379.4]
  wire [7:0] _T_12013; // @[Mux.scala 46:16:@10380.4]
  wire  _T_12014; // @[Mux.scala 46:19:@10381.4]
  wire [7:0] _T_12015; // @[Mux.scala 46:16:@10382.4]
  wire  _T_12016; // @[Mux.scala 46:19:@10383.4]
  wire [7:0] _T_12017; // @[Mux.scala 46:16:@10384.4]
  wire  _T_12018; // @[Mux.scala 46:19:@10385.4]
  wire [7:0] _T_12019; // @[Mux.scala 46:16:@10386.4]
  wire  _T_12020; // @[Mux.scala 46:19:@10387.4]
  wire [7:0] _T_12021; // @[Mux.scala 46:16:@10388.4]
  wire  _T_12022; // @[Mux.scala 46:19:@10389.4]
  wire [7:0] _T_12023; // @[Mux.scala 46:16:@10390.4]
  wire  _T_12024; // @[Mux.scala 46:19:@10391.4]
  wire [7:0] _T_12025; // @[Mux.scala 46:16:@10392.4]
  wire  _T_12060; // @[Mux.scala 46:19:@10394.4]
  wire [7:0] _T_12061; // @[Mux.scala 46:16:@10395.4]
  wire  _T_12062; // @[Mux.scala 46:19:@10396.4]
  wire [7:0] _T_12063; // @[Mux.scala 46:16:@10397.4]
  wire  _T_12064; // @[Mux.scala 46:19:@10398.4]
  wire [7:0] _T_12065; // @[Mux.scala 46:16:@10399.4]
  wire  _T_12066; // @[Mux.scala 46:19:@10400.4]
  wire [7:0] _T_12067; // @[Mux.scala 46:16:@10401.4]
  wire  _T_12068; // @[Mux.scala 46:19:@10402.4]
  wire [7:0] _T_12069; // @[Mux.scala 46:16:@10403.4]
  wire  _T_12070; // @[Mux.scala 46:19:@10404.4]
  wire [7:0] _T_12071; // @[Mux.scala 46:16:@10405.4]
  wire  _T_12072; // @[Mux.scala 46:19:@10406.4]
  wire [7:0] _T_12073; // @[Mux.scala 46:16:@10407.4]
  wire  _T_12074; // @[Mux.scala 46:19:@10408.4]
  wire [7:0] _T_12075; // @[Mux.scala 46:16:@10409.4]
  wire  _T_12076; // @[Mux.scala 46:19:@10410.4]
  wire [7:0] _T_12077; // @[Mux.scala 46:16:@10411.4]
  wire  _T_12078; // @[Mux.scala 46:19:@10412.4]
  wire [7:0] _T_12079; // @[Mux.scala 46:16:@10413.4]
  wire  _T_12080; // @[Mux.scala 46:19:@10414.4]
  wire [7:0] _T_12081; // @[Mux.scala 46:16:@10415.4]
  wire  _T_12082; // @[Mux.scala 46:19:@10416.4]
  wire [7:0] _T_12083; // @[Mux.scala 46:16:@10417.4]
  wire  _T_12084; // @[Mux.scala 46:19:@10418.4]
  wire [7:0] _T_12085; // @[Mux.scala 46:16:@10419.4]
  wire  _T_12086; // @[Mux.scala 46:19:@10420.4]
  wire [7:0] _T_12087; // @[Mux.scala 46:16:@10421.4]
  wire  _T_12088; // @[Mux.scala 46:19:@10422.4]
  wire [7:0] _T_12089; // @[Mux.scala 46:16:@10423.4]
  wire  _T_12090; // @[Mux.scala 46:19:@10424.4]
  wire [7:0] _T_12091; // @[Mux.scala 46:16:@10425.4]
  wire  _T_12092; // @[Mux.scala 46:19:@10426.4]
  wire [7:0] _T_12093; // @[Mux.scala 46:16:@10427.4]
  wire  _T_12094; // @[Mux.scala 46:19:@10428.4]
  wire [7:0] _T_12095; // @[Mux.scala 46:16:@10429.4]
  wire  _T_12096; // @[Mux.scala 46:19:@10430.4]
  wire [7:0] _T_12097; // @[Mux.scala 46:16:@10431.4]
  wire  _T_12098; // @[Mux.scala 46:19:@10432.4]
  wire [7:0] _T_12099; // @[Mux.scala 46:16:@10433.4]
  wire  _T_12100; // @[Mux.scala 46:19:@10434.4]
  wire [7:0] _T_12101; // @[Mux.scala 46:16:@10435.4]
  wire  _T_12102; // @[Mux.scala 46:19:@10436.4]
  wire [7:0] _T_12103; // @[Mux.scala 46:16:@10437.4]
  wire  _T_12104; // @[Mux.scala 46:19:@10438.4]
  wire [7:0] _T_12105; // @[Mux.scala 46:16:@10439.4]
  wire  _T_12106; // @[Mux.scala 46:19:@10440.4]
  wire [7:0] _T_12107; // @[Mux.scala 46:16:@10441.4]
  wire  _T_12108; // @[Mux.scala 46:19:@10442.4]
  wire [7:0] _T_12109; // @[Mux.scala 46:16:@10443.4]
  wire  _T_12110; // @[Mux.scala 46:19:@10444.4]
  wire [7:0] _T_12111; // @[Mux.scala 46:16:@10445.4]
  wire  _T_12112; // @[Mux.scala 46:19:@10446.4]
  wire [7:0] _T_12113; // @[Mux.scala 46:16:@10447.4]
  wire  _T_12114; // @[Mux.scala 46:19:@10448.4]
  wire [7:0] _T_12115; // @[Mux.scala 46:16:@10449.4]
  wire  _T_12116; // @[Mux.scala 46:19:@10450.4]
  wire [7:0] _T_12117; // @[Mux.scala 46:16:@10451.4]
  wire  _T_12118; // @[Mux.scala 46:19:@10452.4]
  wire [7:0] _T_12119; // @[Mux.scala 46:16:@10453.4]
  wire  _T_12120; // @[Mux.scala 46:19:@10454.4]
  wire [7:0] _T_12121; // @[Mux.scala 46:16:@10455.4]
  wire  _T_12122; // @[Mux.scala 46:19:@10456.4]
  wire [7:0] _T_12123; // @[Mux.scala 46:16:@10457.4]
  wire  _T_12124; // @[Mux.scala 46:19:@10458.4]
  wire [7:0] _T_12125; // @[Mux.scala 46:16:@10459.4]
  wire  _T_12161; // @[Mux.scala 46:19:@10461.4]
  wire [7:0] _T_12162; // @[Mux.scala 46:16:@10462.4]
  wire  _T_12163; // @[Mux.scala 46:19:@10463.4]
  wire [7:0] _T_12164; // @[Mux.scala 46:16:@10464.4]
  wire  _T_12165; // @[Mux.scala 46:19:@10465.4]
  wire [7:0] _T_12166; // @[Mux.scala 46:16:@10466.4]
  wire  _T_12167; // @[Mux.scala 46:19:@10467.4]
  wire [7:0] _T_12168; // @[Mux.scala 46:16:@10468.4]
  wire  _T_12169; // @[Mux.scala 46:19:@10469.4]
  wire [7:0] _T_12170; // @[Mux.scala 46:16:@10470.4]
  wire  _T_12171; // @[Mux.scala 46:19:@10471.4]
  wire [7:0] _T_12172; // @[Mux.scala 46:16:@10472.4]
  wire  _T_12173; // @[Mux.scala 46:19:@10473.4]
  wire [7:0] _T_12174; // @[Mux.scala 46:16:@10474.4]
  wire  _T_12175; // @[Mux.scala 46:19:@10475.4]
  wire [7:0] _T_12176; // @[Mux.scala 46:16:@10476.4]
  wire  _T_12177; // @[Mux.scala 46:19:@10477.4]
  wire [7:0] _T_12178; // @[Mux.scala 46:16:@10478.4]
  wire  _T_12179; // @[Mux.scala 46:19:@10479.4]
  wire [7:0] _T_12180; // @[Mux.scala 46:16:@10480.4]
  wire  _T_12181; // @[Mux.scala 46:19:@10481.4]
  wire [7:0] _T_12182; // @[Mux.scala 46:16:@10482.4]
  wire  _T_12183; // @[Mux.scala 46:19:@10483.4]
  wire [7:0] _T_12184; // @[Mux.scala 46:16:@10484.4]
  wire  _T_12185; // @[Mux.scala 46:19:@10485.4]
  wire [7:0] _T_12186; // @[Mux.scala 46:16:@10486.4]
  wire  _T_12187; // @[Mux.scala 46:19:@10487.4]
  wire [7:0] _T_12188; // @[Mux.scala 46:16:@10488.4]
  wire  _T_12189; // @[Mux.scala 46:19:@10489.4]
  wire [7:0] _T_12190; // @[Mux.scala 46:16:@10490.4]
  wire  _T_12191; // @[Mux.scala 46:19:@10491.4]
  wire [7:0] _T_12192; // @[Mux.scala 46:16:@10492.4]
  wire  _T_12193; // @[Mux.scala 46:19:@10493.4]
  wire [7:0] _T_12194; // @[Mux.scala 46:16:@10494.4]
  wire  _T_12195; // @[Mux.scala 46:19:@10495.4]
  wire [7:0] _T_12196; // @[Mux.scala 46:16:@10496.4]
  wire  _T_12197; // @[Mux.scala 46:19:@10497.4]
  wire [7:0] _T_12198; // @[Mux.scala 46:16:@10498.4]
  wire  _T_12199; // @[Mux.scala 46:19:@10499.4]
  wire [7:0] _T_12200; // @[Mux.scala 46:16:@10500.4]
  wire  _T_12201; // @[Mux.scala 46:19:@10501.4]
  wire [7:0] _T_12202; // @[Mux.scala 46:16:@10502.4]
  wire  _T_12203; // @[Mux.scala 46:19:@10503.4]
  wire [7:0] _T_12204; // @[Mux.scala 46:16:@10504.4]
  wire  _T_12205; // @[Mux.scala 46:19:@10505.4]
  wire [7:0] _T_12206; // @[Mux.scala 46:16:@10506.4]
  wire  _T_12207; // @[Mux.scala 46:19:@10507.4]
  wire [7:0] _T_12208; // @[Mux.scala 46:16:@10508.4]
  wire  _T_12209; // @[Mux.scala 46:19:@10509.4]
  wire [7:0] _T_12210; // @[Mux.scala 46:16:@10510.4]
  wire  _T_12211; // @[Mux.scala 46:19:@10511.4]
  wire [7:0] _T_12212; // @[Mux.scala 46:16:@10512.4]
  wire  _T_12213; // @[Mux.scala 46:19:@10513.4]
  wire [7:0] _T_12214; // @[Mux.scala 46:16:@10514.4]
  wire  _T_12215; // @[Mux.scala 46:19:@10515.4]
  wire [7:0] _T_12216; // @[Mux.scala 46:16:@10516.4]
  wire  _T_12217; // @[Mux.scala 46:19:@10517.4]
  wire [7:0] _T_12218; // @[Mux.scala 46:16:@10518.4]
  wire  _T_12219; // @[Mux.scala 46:19:@10519.4]
  wire [7:0] _T_12220; // @[Mux.scala 46:16:@10520.4]
  wire  _T_12221; // @[Mux.scala 46:19:@10521.4]
  wire [7:0] _T_12222; // @[Mux.scala 46:16:@10522.4]
  wire  _T_12223; // @[Mux.scala 46:19:@10523.4]
  wire [7:0] _T_12224; // @[Mux.scala 46:16:@10524.4]
  wire  _T_12225; // @[Mux.scala 46:19:@10525.4]
  wire [7:0] _T_12226; // @[Mux.scala 46:16:@10526.4]
  wire  _T_12227; // @[Mux.scala 46:19:@10527.4]
  wire [7:0] _T_12228; // @[Mux.scala 46:16:@10528.4]
  wire  _T_12265; // @[Mux.scala 46:19:@10530.4]
  wire [7:0] _T_12266; // @[Mux.scala 46:16:@10531.4]
  wire  _T_12267; // @[Mux.scala 46:19:@10532.4]
  wire [7:0] _T_12268; // @[Mux.scala 46:16:@10533.4]
  wire  _T_12269; // @[Mux.scala 46:19:@10534.4]
  wire [7:0] _T_12270; // @[Mux.scala 46:16:@10535.4]
  wire  _T_12271; // @[Mux.scala 46:19:@10536.4]
  wire [7:0] _T_12272; // @[Mux.scala 46:16:@10537.4]
  wire  _T_12273; // @[Mux.scala 46:19:@10538.4]
  wire [7:0] _T_12274; // @[Mux.scala 46:16:@10539.4]
  wire  _T_12275; // @[Mux.scala 46:19:@10540.4]
  wire [7:0] _T_12276; // @[Mux.scala 46:16:@10541.4]
  wire  _T_12277; // @[Mux.scala 46:19:@10542.4]
  wire [7:0] _T_12278; // @[Mux.scala 46:16:@10543.4]
  wire  _T_12279; // @[Mux.scala 46:19:@10544.4]
  wire [7:0] _T_12280; // @[Mux.scala 46:16:@10545.4]
  wire  _T_12281; // @[Mux.scala 46:19:@10546.4]
  wire [7:0] _T_12282; // @[Mux.scala 46:16:@10547.4]
  wire  _T_12283; // @[Mux.scala 46:19:@10548.4]
  wire [7:0] _T_12284; // @[Mux.scala 46:16:@10549.4]
  wire  _T_12285; // @[Mux.scala 46:19:@10550.4]
  wire [7:0] _T_12286; // @[Mux.scala 46:16:@10551.4]
  wire  _T_12287; // @[Mux.scala 46:19:@10552.4]
  wire [7:0] _T_12288; // @[Mux.scala 46:16:@10553.4]
  wire  _T_12289; // @[Mux.scala 46:19:@10554.4]
  wire [7:0] _T_12290; // @[Mux.scala 46:16:@10555.4]
  wire  _T_12291; // @[Mux.scala 46:19:@10556.4]
  wire [7:0] _T_12292; // @[Mux.scala 46:16:@10557.4]
  wire  _T_12293; // @[Mux.scala 46:19:@10558.4]
  wire [7:0] _T_12294; // @[Mux.scala 46:16:@10559.4]
  wire  _T_12295; // @[Mux.scala 46:19:@10560.4]
  wire [7:0] _T_12296; // @[Mux.scala 46:16:@10561.4]
  wire  _T_12297; // @[Mux.scala 46:19:@10562.4]
  wire [7:0] _T_12298; // @[Mux.scala 46:16:@10563.4]
  wire  _T_12299; // @[Mux.scala 46:19:@10564.4]
  wire [7:0] _T_12300; // @[Mux.scala 46:16:@10565.4]
  wire  _T_12301; // @[Mux.scala 46:19:@10566.4]
  wire [7:0] _T_12302; // @[Mux.scala 46:16:@10567.4]
  wire  _T_12303; // @[Mux.scala 46:19:@10568.4]
  wire [7:0] _T_12304; // @[Mux.scala 46:16:@10569.4]
  wire  _T_12305; // @[Mux.scala 46:19:@10570.4]
  wire [7:0] _T_12306; // @[Mux.scala 46:16:@10571.4]
  wire  _T_12307; // @[Mux.scala 46:19:@10572.4]
  wire [7:0] _T_12308; // @[Mux.scala 46:16:@10573.4]
  wire  _T_12309; // @[Mux.scala 46:19:@10574.4]
  wire [7:0] _T_12310; // @[Mux.scala 46:16:@10575.4]
  wire  _T_12311; // @[Mux.scala 46:19:@10576.4]
  wire [7:0] _T_12312; // @[Mux.scala 46:16:@10577.4]
  wire  _T_12313; // @[Mux.scala 46:19:@10578.4]
  wire [7:0] _T_12314; // @[Mux.scala 46:16:@10579.4]
  wire  _T_12315; // @[Mux.scala 46:19:@10580.4]
  wire [7:0] _T_12316; // @[Mux.scala 46:16:@10581.4]
  wire  _T_12317; // @[Mux.scala 46:19:@10582.4]
  wire [7:0] _T_12318; // @[Mux.scala 46:16:@10583.4]
  wire  _T_12319; // @[Mux.scala 46:19:@10584.4]
  wire [7:0] _T_12320; // @[Mux.scala 46:16:@10585.4]
  wire  _T_12321; // @[Mux.scala 46:19:@10586.4]
  wire [7:0] _T_12322; // @[Mux.scala 46:16:@10587.4]
  wire  _T_12323; // @[Mux.scala 46:19:@10588.4]
  wire [7:0] _T_12324; // @[Mux.scala 46:16:@10589.4]
  wire  _T_12325; // @[Mux.scala 46:19:@10590.4]
  wire [7:0] _T_12326; // @[Mux.scala 46:16:@10591.4]
  wire  _T_12327; // @[Mux.scala 46:19:@10592.4]
  wire [7:0] _T_12328; // @[Mux.scala 46:16:@10593.4]
  wire  _T_12329; // @[Mux.scala 46:19:@10594.4]
  wire [7:0] _T_12330; // @[Mux.scala 46:16:@10595.4]
  wire  _T_12331; // @[Mux.scala 46:19:@10596.4]
  wire [7:0] _T_12332; // @[Mux.scala 46:16:@10597.4]
  wire  _T_12333; // @[Mux.scala 46:19:@10598.4]
  wire [7:0] _T_12334; // @[Mux.scala 46:16:@10599.4]
  wire  _T_12372; // @[Mux.scala 46:19:@10601.4]
  wire [7:0] _T_12373; // @[Mux.scala 46:16:@10602.4]
  wire  _T_12374; // @[Mux.scala 46:19:@10603.4]
  wire [7:0] _T_12375; // @[Mux.scala 46:16:@10604.4]
  wire  _T_12376; // @[Mux.scala 46:19:@10605.4]
  wire [7:0] _T_12377; // @[Mux.scala 46:16:@10606.4]
  wire  _T_12378; // @[Mux.scala 46:19:@10607.4]
  wire [7:0] _T_12379; // @[Mux.scala 46:16:@10608.4]
  wire  _T_12380; // @[Mux.scala 46:19:@10609.4]
  wire [7:0] _T_12381; // @[Mux.scala 46:16:@10610.4]
  wire  _T_12382; // @[Mux.scala 46:19:@10611.4]
  wire [7:0] _T_12383; // @[Mux.scala 46:16:@10612.4]
  wire  _T_12384; // @[Mux.scala 46:19:@10613.4]
  wire [7:0] _T_12385; // @[Mux.scala 46:16:@10614.4]
  wire  _T_12386; // @[Mux.scala 46:19:@10615.4]
  wire [7:0] _T_12387; // @[Mux.scala 46:16:@10616.4]
  wire  _T_12388; // @[Mux.scala 46:19:@10617.4]
  wire [7:0] _T_12389; // @[Mux.scala 46:16:@10618.4]
  wire  _T_12390; // @[Mux.scala 46:19:@10619.4]
  wire [7:0] _T_12391; // @[Mux.scala 46:16:@10620.4]
  wire  _T_12392; // @[Mux.scala 46:19:@10621.4]
  wire [7:0] _T_12393; // @[Mux.scala 46:16:@10622.4]
  wire  _T_12394; // @[Mux.scala 46:19:@10623.4]
  wire [7:0] _T_12395; // @[Mux.scala 46:16:@10624.4]
  wire  _T_12396; // @[Mux.scala 46:19:@10625.4]
  wire [7:0] _T_12397; // @[Mux.scala 46:16:@10626.4]
  wire  _T_12398; // @[Mux.scala 46:19:@10627.4]
  wire [7:0] _T_12399; // @[Mux.scala 46:16:@10628.4]
  wire  _T_12400; // @[Mux.scala 46:19:@10629.4]
  wire [7:0] _T_12401; // @[Mux.scala 46:16:@10630.4]
  wire  _T_12402; // @[Mux.scala 46:19:@10631.4]
  wire [7:0] _T_12403; // @[Mux.scala 46:16:@10632.4]
  wire  _T_12404; // @[Mux.scala 46:19:@10633.4]
  wire [7:0] _T_12405; // @[Mux.scala 46:16:@10634.4]
  wire  _T_12406; // @[Mux.scala 46:19:@10635.4]
  wire [7:0] _T_12407; // @[Mux.scala 46:16:@10636.4]
  wire  _T_12408; // @[Mux.scala 46:19:@10637.4]
  wire [7:0] _T_12409; // @[Mux.scala 46:16:@10638.4]
  wire  _T_12410; // @[Mux.scala 46:19:@10639.4]
  wire [7:0] _T_12411; // @[Mux.scala 46:16:@10640.4]
  wire  _T_12412; // @[Mux.scala 46:19:@10641.4]
  wire [7:0] _T_12413; // @[Mux.scala 46:16:@10642.4]
  wire  _T_12414; // @[Mux.scala 46:19:@10643.4]
  wire [7:0] _T_12415; // @[Mux.scala 46:16:@10644.4]
  wire  _T_12416; // @[Mux.scala 46:19:@10645.4]
  wire [7:0] _T_12417; // @[Mux.scala 46:16:@10646.4]
  wire  _T_12418; // @[Mux.scala 46:19:@10647.4]
  wire [7:0] _T_12419; // @[Mux.scala 46:16:@10648.4]
  wire  _T_12420; // @[Mux.scala 46:19:@10649.4]
  wire [7:0] _T_12421; // @[Mux.scala 46:16:@10650.4]
  wire  _T_12422; // @[Mux.scala 46:19:@10651.4]
  wire [7:0] _T_12423; // @[Mux.scala 46:16:@10652.4]
  wire  _T_12424; // @[Mux.scala 46:19:@10653.4]
  wire [7:0] _T_12425; // @[Mux.scala 46:16:@10654.4]
  wire  _T_12426; // @[Mux.scala 46:19:@10655.4]
  wire [7:0] _T_12427; // @[Mux.scala 46:16:@10656.4]
  wire  _T_12428; // @[Mux.scala 46:19:@10657.4]
  wire [7:0] _T_12429; // @[Mux.scala 46:16:@10658.4]
  wire  _T_12430; // @[Mux.scala 46:19:@10659.4]
  wire [7:0] _T_12431; // @[Mux.scala 46:16:@10660.4]
  wire  _T_12432; // @[Mux.scala 46:19:@10661.4]
  wire [7:0] _T_12433; // @[Mux.scala 46:16:@10662.4]
  wire  _T_12434; // @[Mux.scala 46:19:@10663.4]
  wire [7:0] _T_12435; // @[Mux.scala 46:16:@10664.4]
  wire  _T_12436; // @[Mux.scala 46:19:@10665.4]
  wire [7:0] _T_12437; // @[Mux.scala 46:16:@10666.4]
  wire  _T_12438; // @[Mux.scala 46:19:@10667.4]
  wire [7:0] _T_12439; // @[Mux.scala 46:16:@10668.4]
  wire  _T_12440; // @[Mux.scala 46:19:@10669.4]
  wire [7:0] _T_12441; // @[Mux.scala 46:16:@10670.4]
  wire  _T_12442; // @[Mux.scala 46:19:@10671.4]
  wire [7:0] _T_12443; // @[Mux.scala 46:16:@10672.4]
  wire  _T_12482; // @[Mux.scala 46:19:@10674.4]
  wire [7:0] _T_12483; // @[Mux.scala 46:16:@10675.4]
  wire  _T_12484; // @[Mux.scala 46:19:@10676.4]
  wire [7:0] _T_12485; // @[Mux.scala 46:16:@10677.4]
  wire  _T_12486; // @[Mux.scala 46:19:@10678.4]
  wire [7:0] _T_12487; // @[Mux.scala 46:16:@10679.4]
  wire  _T_12488; // @[Mux.scala 46:19:@10680.4]
  wire [7:0] _T_12489; // @[Mux.scala 46:16:@10681.4]
  wire  _T_12490; // @[Mux.scala 46:19:@10682.4]
  wire [7:0] _T_12491; // @[Mux.scala 46:16:@10683.4]
  wire  _T_12492; // @[Mux.scala 46:19:@10684.4]
  wire [7:0] _T_12493; // @[Mux.scala 46:16:@10685.4]
  wire  _T_12494; // @[Mux.scala 46:19:@10686.4]
  wire [7:0] _T_12495; // @[Mux.scala 46:16:@10687.4]
  wire  _T_12496; // @[Mux.scala 46:19:@10688.4]
  wire [7:0] _T_12497; // @[Mux.scala 46:16:@10689.4]
  wire  _T_12498; // @[Mux.scala 46:19:@10690.4]
  wire [7:0] _T_12499; // @[Mux.scala 46:16:@10691.4]
  wire  _T_12500; // @[Mux.scala 46:19:@10692.4]
  wire [7:0] _T_12501; // @[Mux.scala 46:16:@10693.4]
  wire  _T_12502; // @[Mux.scala 46:19:@10694.4]
  wire [7:0] _T_12503; // @[Mux.scala 46:16:@10695.4]
  wire  _T_12504; // @[Mux.scala 46:19:@10696.4]
  wire [7:0] _T_12505; // @[Mux.scala 46:16:@10697.4]
  wire  _T_12506; // @[Mux.scala 46:19:@10698.4]
  wire [7:0] _T_12507; // @[Mux.scala 46:16:@10699.4]
  wire  _T_12508; // @[Mux.scala 46:19:@10700.4]
  wire [7:0] _T_12509; // @[Mux.scala 46:16:@10701.4]
  wire  _T_12510; // @[Mux.scala 46:19:@10702.4]
  wire [7:0] _T_12511; // @[Mux.scala 46:16:@10703.4]
  wire  _T_12512; // @[Mux.scala 46:19:@10704.4]
  wire [7:0] _T_12513; // @[Mux.scala 46:16:@10705.4]
  wire  _T_12514; // @[Mux.scala 46:19:@10706.4]
  wire [7:0] _T_12515; // @[Mux.scala 46:16:@10707.4]
  wire  _T_12516; // @[Mux.scala 46:19:@10708.4]
  wire [7:0] _T_12517; // @[Mux.scala 46:16:@10709.4]
  wire  _T_12518; // @[Mux.scala 46:19:@10710.4]
  wire [7:0] _T_12519; // @[Mux.scala 46:16:@10711.4]
  wire  _T_12520; // @[Mux.scala 46:19:@10712.4]
  wire [7:0] _T_12521; // @[Mux.scala 46:16:@10713.4]
  wire  _T_12522; // @[Mux.scala 46:19:@10714.4]
  wire [7:0] _T_12523; // @[Mux.scala 46:16:@10715.4]
  wire  _T_12524; // @[Mux.scala 46:19:@10716.4]
  wire [7:0] _T_12525; // @[Mux.scala 46:16:@10717.4]
  wire  _T_12526; // @[Mux.scala 46:19:@10718.4]
  wire [7:0] _T_12527; // @[Mux.scala 46:16:@10719.4]
  wire  _T_12528; // @[Mux.scala 46:19:@10720.4]
  wire [7:0] _T_12529; // @[Mux.scala 46:16:@10721.4]
  wire  _T_12530; // @[Mux.scala 46:19:@10722.4]
  wire [7:0] _T_12531; // @[Mux.scala 46:16:@10723.4]
  wire  _T_12532; // @[Mux.scala 46:19:@10724.4]
  wire [7:0] _T_12533; // @[Mux.scala 46:16:@10725.4]
  wire  _T_12534; // @[Mux.scala 46:19:@10726.4]
  wire [7:0] _T_12535; // @[Mux.scala 46:16:@10727.4]
  wire  _T_12536; // @[Mux.scala 46:19:@10728.4]
  wire [7:0] _T_12537; // @[Mux.scala 46:16:@10729.4]
  wire  _T_12538; // @[Mux.scala 46:19:@10730.4]
  wire [7:0] _T_12539; // @[Mux.scala 46:16:@10731.4]
  wire  _T_12540; // @[Mux.scala 46:19:@10732.4]
  wire [7:0] _T_12541; // @[Mux.scala 46:16:@10733.4]
  wire  _T_12542; // @[Mux.scala 46:19:@10734.4]
  wire [7:0] _T_12543; // @[Mux.scala 46:16:@10735.4]
  wire  _T_12544; // @[Mux.scala 46:19:@10736.4]
  wire [7:0] _T_12545; // @[Mux.scala 46:16:@10737.4]
  wire  _T_12546; // @[Mux.scala 46:19:@10738.4]
  wire [7:0] _T_12547; // @[Mux.scala 46:16:@10739.4]
  wire  _T_12548; // @[Mux.scala 46:19:@10740.4]
  wire [7:0] _T_12549; // @[Mux.scala 46:16:@10741.4]
  wire  _T_12550; // @[Mux.scala 46:19:@10742.4]
  wire [7:0] _T_12551; // @[Mux.scala 46:16:@10743.4]
  wire  _T_12552; // @[Mux.scala 46:19:@10744.4]
  wire [7:0] _T_12553; // @[Mux.scala 46:16:@10745.4]
  wire  _T_12554; // @[Mux.scala 46:19:@10746.4]
  wire [7:0] _T_12555; // @[Mux.scala 46:16:@10747.4]
  wire  _T_12595; // @[Mux.scala 46:19:@10749.4]
  wire [7:0] _T_12596; // @[Mux.scala 46:16:@10750.4]
  wire  _T_12597; // @[Mux.scala 46:19:@10751.4]
  wire [7:0] _T_12598; // @[Mux.scala 46:16:@10752.4]
  wire  _T_12599; // @[Mux.scala 46:19:@10753.4]
  wire [7:0] _T_12600; // @[Mux.scala 46:16:@10754.4]
  wire  _T_12601; // @[Mux.scala 46:19:@10755.4]
  wire [7:0] _T_12602; // @[Mux.scala 46:16:@10756.4]
  wire  _T_12603; // @[Mux.scala 46:19:@10757.4]
  wire [7:0] _T_12604; // @[Mux.scala 46:16:@10758.4]
  wire  _T_12605; // @[Mux.scala 46:19:@10759.4]
  wire [7:0] _T_12606; // @[Mux.scala 46:16:@10760.4]
  wire  _T_12607; // @[Mux.scala 46:19:@10761.4]
  wire [7:0] _T_12608; // @[Mux.scala 46:16:@10762.4]
  wire  _T_12609; // @[Mux.scala 46:19:@10763.4]
  wire [7:0] _T_12610; // @[Mux.scala 46:16:@10764.4]
  wire  _T_12611; // @[Mux.scala 46:19:@10765.4]
  wire [7:0] _T_12612; // @[Mux.scala 46:16:@10766.4]
  wire  _T_12613; // @[Mux.scala 46:19:@10767.4]
  wire [7:0] _T_12614; // @[Mux.scala 46:16:@10768.4]
  wire  _T_12615; // @[Mux.scala 46:19:@10769.4]
  wire [7:0] _T_12616; // @[Mux.scala 46:16:@10770.4]
  wire  _T_12617; // @[Mux.scala 46:19:@10771.4]
  wire [7:0] _T_12618; // @[Mux.scala 46:16:@10772.4]
  wire  _T_12619; // @[Mux.scala 46:19:@10773.4]
  wire [7:0] _T_12620; // @[Mux.scala 46:16:@10774.4]
  wire  _T_12621; // @[Mux.scala 46:19:@10775.4]
  wire [7:0] _T_12622; // @[Mux.scala 46:16:@10776.4]
  wire  _T_12623; // @[Mux.scala 46:19:@10777.4]
  wire [7:0] _T_12624; // @[Mux.scala 46:16:@10778.4]
  wire  _T_12625; // @[Mux.scala 46:19:@10779.4]
  wire [7:0] _T_12626; // @[Mux.scala 46:16:@10780.4]
  wire  _T_12627; // @[Mux.scala 46:19:@10781.4]
  wire [7:0] _T_12628; // @[Mux.scala 46:16:@10782.4]
  wire  _T_12629; // @[Mux.scala 46:19:@10783.4]
  wire [7:0] _T_12630; // @[Mux.scala 46:16:@10784.4]
  wire  _T_12631; // @[Mux.scala 46:19:@10785.4]
  wire [7:0] _T_12632; // @[Mux.scala 46:16:@10786.4]
  wire  _T_12633; // @[Mux.scala 46:19:@10787.4]
  wire [7:0] _T_12634; // @[Mux.scala 46:16:@10788.4]
  wire  _T_12635; // @[Mux.scala 46:19:@10789.4]
  wire [7:0] _T_12636; // @[Mux.scala 46:16:@10790.4]
  wire  _T_12637; // @[Mux.scala 46:19:@10791.4]
  wire [7:0] _T_12638; // @[Mux.scala 46:16:@10792.4]
  wire  _T_12639; // @[Mux.scala 46:19:@10793.4]
  wire [7:0] _T_12640; // @[Mux.scala 46:16:@10794.4]
  wire  _T_12641; // @[Mux.scala 46:19:@10795.4]
  wire [7:0] _T_12642; // @[Mux.scala 46:16:@10796.4]
  wire  _T_12643; // @[Mux.scala 46:19:@10797.4]
  wire [7:0] _T_12644; // @[Mux.scala 46:16:@10798.4]
  wire  _T_12645; // @[Mux.scala 46:19:@10799.4]
  wire [7:0] _T_12646; // @[Mux.scala 46:16:@10800.4]
  wire  _T_12647; // @[Mux.scala 46:19:@10801.4]
  wire [7:0] _T_12648; // @[Mux.scala 46:16:@10802.4]
  wire  _T_12649; // @[Mux.scala 46:19:@10803.4]
  wire [7:0] _T_12650; // @[Mux.scala 46:16:@10804.4]
  wire  _T_12651; // @[Mux.scala 46:19:@10805.4]
  wire [7:0] _T_12652; // @[Mux.scala 46:16:@10806.4]
  wire  _T_12653; // @[Mux.scala 46:19:@10807.4]
  wire [7:0] _T_12654; // @[Mux.scala 46:16:@10808.4]
  wire  _T_12655; // @[Mux.scala 46:19:@10809.4]
  wire [7:0] _T_12656; // @[Mux.scala 46:16:@10810.4]
  wire  _T_12657; // @[Mux.scala 46:19:@10811.4]
  wire [7:0] _T_12658; // @[Mux.scala 46:16:@10812.4]
  wire  _T_12659; // @[Mux.scala 46:19:@10813.4]
  wire [7:0] _T_12660; // @[Mux.scala 46:16:@10814.4]
  wire  _T_12661; // @[Mux.scala 46:19:@10815.4]
  wire [7:0] _T_12662; // @[Mux.scala 46:16:@10816.4]
  wire  _T_12663; // @[Mux.scala 46:19:@10817.4]
  wire [7:0] _T_12664; // @[Mux.scala 46:16:@10818.4]
  wire  _T_12665; // @[Mux.scala 46:19:@10819.4]
  wire [7:0] _T_12666; // @[Mux.scala 46:16:@10820.4]
  wire  _T_12667; // @[Mux.scala 46:19:@10821.4]
  wire [7:0] _T_12668; // @[Mux.scala 46:16:@10822.4]
  wire  _T_12669; // @[Mux.scala 46:19:@10823.4]
  wire [7:0] _T_12670; // @[Mux.scala 46:16:@10824.4]
  wire  _T_12711; // @[Mux.scala 46:19:@10826.4]
  wire [7:0] _T_12712; // @[Mux.scala 46:16:@10827.4]
  wire  _T_12713; // @[Mux.scala 46:19:@10828.4]
  wire [7:0] _T_12714; // @[Mux.scala 46:16:@10829.4]
  wire  _T_12715; // @[Mux.scala 46:19:@10830.4]
  wire [7:0] _T_12716; // @[Mux.scala 46:16:@10831.4]
  wire  _T_12717; // @[Mux.scala 46:19:@10832.4]
  wire [7:0] _T_12718; // @[Mux.scala 46:16:@10833.4]
  wire  _T_12719; // @[Mux.scala 46:19:@10834.4]
  wire [7:0] _T_12720; // @[Mux.scala 46:16:@10835.4]
  wire  _T_12721; // @[Mux.scala 46:19:@10836.4]
  wire [7:0] _T_12722; // @[Mux.scala 46:16:@10837.4]
  wire  _T_12723; // @[Mux.scala 46:19:@10838.4]
  wire [7:0] _T_12724; // @[Mux.scala 46:16:@10839.4]
  wire  _T_12725; // @[Mux.scala 46:19:@10840.4]
  wire [7:0] _T_12726; // @[Mux.scala 46:16:@10841.4]
  wire  _T_12727; // @[Mux.scala 46:19:@10842.4]
  wire [7:0] _T_12728; // @[Mux.scala 46:16:@10843.4]
  wire  _T_12729; // @[Mux.scala 46:19:@10844.4]
  wire [7:0] _T_12730; // @[Mux.scala 46:16:@10845.4]
  wire  _T_12731; // @[Mux.scala 46:19:@10846.4]
  wire [7:0] _T_12732; // @[Mux.scala 46:16:@10847.4]
  wire  _T_12733; // @[Mux.scala 46:19:@10848.4]
  wire [7:0] _T_12734; // @[Mux.scala 46:16:@10849.4]
  wire  _T_12735; // @[Mux.scala 46:19:@10850.4]
  wire [7:0] _T_12736; // @[Mux.scala 46:16:@10851.4]
  wire  _T_12737; // @[Mux.scala 46:19:@10852.4]
  wire [7:0] _T_12738; // @[Mux.scala 46:16:@10853.4]
  wire  _T_12739; // @[Mux.scala 46:19:@10854.4]
  wire [7:0] _T_12740; // @[Mux.scala 46:16:@10855.4]
  wire  _T_12741; // @[Mux.scala 46:19:@10856.4]
  wire [7:0] _T_12742; // @[Mux.scala 46:16:@10857.4]
  wire  _T_12743; // @[Mux.scala 46:19:@10858.4]
  wire [7:0] _T_12744; // @[Mux.scala 46:16:@10859.4]
  wire  _T_12745; // @[Mux.scala 46:19:@10860.4]
  wire [7:0] _T_12746; // @[Mux.scala 46:16:@10861.4]
  wire  _T_12747; // @[Mux.scala 46:19:@10862.4]
  wire [7:0] _T_12748; // @[Mux.scala 46:16:@10863.4]
  wire  _T_12749; // @[Mux.scala 46:19:@10864.4]
  wire [7:0] _T_12750; // @[Mux.scala 46:16:@10865.4]
  wire  _T_12751; // @[Mux.scala 46:19:@10866.4]
  wire [7:0] _T_12752; // @[Mux.scala 46:16:@10867.4]
  wire  _T_12753; // @[Mux.scala 46:19:@10868.4]
  wire [7:0] _T_12754; // @[Mux.scala 46:16:@10869.4]
  wire  _T_12755; // @[Mux.scala 46:19:@10870.4]
  wire [7:0] _T_12756; // @[Mux.scala 46:16:@10871.4]
  wire  _T_12757; // @[Mux.scala 46:19:@10872.4]
  wire [7:0] _T_12758; // @[Mux.scala 46:16:@10873.4]
  wire  _T_12759; // @[Mux.scala 46:19:@10874.4]
  wire [7:0] _T_12760; // @[Mux.scala 46:16:@10875.4]
  wire  _T_12761; // @[Mux.scala 46:19:@10876.4]
  wire [7:0] _T_12762; // @[Mux.scala 46:16:@10877.4]
  wire  _T_12763; // @[Mux.scala 46:19:@10878.4]
  wire [7:0] _T_12764; // @[Mux.scala 46:16:@10879.4]
  wire  _T_12765; // @[Mux.scala 46:19:@10880.4]
  wire [7:0] _T_12766; // @[Mux.scala 46:16:@10881.4]
  wire  _T_12767; // @[Mux.scala 46:19:@10882.4]
  wire [7:0] _T_12768; // @[Mux.scala 46:16:@10883.4]
  wire  _T_12769; // @[Mux.scala 46:19:@10884.4]
  wire [7:0] _T_12770; // @[Mux.scala 46:16:@10885.4]
  wire  _T_12771; // @[Mux.scala 46:19:@10886.4]
  wire [7:0] _T_12772; // @[Mux.scala 46:16:@10887.4]
  wire  _T_12773; // @[Mux.scala 46:19:@10888.4]
  wire [7:0] _T_12774; // @[Mux.scala 46:16:@10889.4]
  wire  _T_12775; // @[Mux.scala 46:19:@10890.4]
  wire [7:0] _T_12776; // @[Mux.scala 46:16:@10891.4]
  wire  _T_12777; // @[Mux.scala 46:19:@10892.4]
  wire [7:0] _T_12778; // @[Mux.scala 46:16:@10893.4]
  wire  _T_12779; // @[Mux.scala 46:19:@10894.4]
  wire [7:0] _T_12780; // @[Mux.scala 46:16:@10895.4]
  wire  _T_12781; // @[Mux.scala 46:19:@10896.4]
  wire [7:0] _T_12782; // @[Mux.scala 46:16:@10897.4]
  wire  _T_12783; // @[Mux.scala 46:19:@10898.4]
  wire [7:0] _T_12784; // @[Mux.scala 46:16:@10899.4]
  wire  _T_12785; // @[Mux.scala 46:19:@10900.4]
  wire [7:0] _T_12786; // @[Mux.scala 46:16:@10901.4]
  wire  _T_12787; // @[Mux.scala 46:19:@10902.4]
  wire [7:0] _T_12788; // @[Mux.scala 46:16:@10903.4]
  wire  _T_12830; // @[Mux.scala 46:19:@10905.4]
  wire [7:0] _T_12831; // @[Mux.scala 46:16:@10906.4]
  wire  _T_12832; // @[Mux.scala 46:19:@10907.4]
  wire [7:0] _T_12833; // @[Mux.scala 46:16:@10908.4]
  wire  _T_12834; // @[Mux.scala 46:19:@10909.4]
  wire [7:0] _T_12835; // @[Mux.scala 46:16:@10910.4]
  wire  _T_12836; // @[Mux.scala 46:19:@10911.4]
  wire [7:0] _T_12837; // @[Mux.scala 46:16:@10912.4]
  wire  _T_12838; // @[Mux.scala 46:19:@10913.4]
  wire [7:0] _T_12839; // @[Mux.scala 46:16:@10914.4]
  wire  _T_12840; // @[Mux.scala 46:19:@10915.4]
  wire [7:0] _T_12841; // @[Mux.scala 46:16:@10916.4]
  wire  _T_12842; // @[Mux.scala 46:19:@10917.4]
  wire [7:0] _T_12843; // @[Mux.scala 46:16:@10918.4]
  wire  _T_12844; // @[Mux.scala 46:19:@10919.4]
  wire [7:0] _T_12845; // @[Mux.scala 46:16:@10920.4]
  wire  _T_12846; // @[Mux.scala 46:19:@10921.4]
  wire [7:0] _T_12847; // @[Mux.scala 46:16:@10922.4]
  wire  _T_12848; // @[Mux.scala 46:19:@10923.4]
  wire [7:0] _T_12849; // @[Mux.scala 46:16:@10924.4]
  wire  _T_12850; // @[Mux.scala 46:19:@10925.4]
  wire [7:0] _T_12851; // @[Mux.scala 46:16:@10926.4]
  wire  _T_12852; // @[Mux.scala 46:19:@10927.4]
  wire [7:0] _T_12853; // @[Mux.scala 46:16:@10928.4]
  wire  _T_12854; // @[Mux.scala 46:19:@10929.4]
  wire [7:0] _T_12855; // @[Mux.scala 46:16:@10930.4]
  wire  _T_12856; // @[Mux.scala 46:19:@10931.4]
  wire [7:0] _T_12857; // @[Mux.scala 46:16:@10932.4]
  wire  _T_12858; // @[Mux.scala 46:19:@10933.4]
  wire [7:0] _T_12859; // @[Mux.scala 46:16:@10934.4]
  wire  _T_12860; // @[Mux.scala 46:19:@10935.4]
  wire [7:0] _T_12861; // @[Mux.scala 46:16:@10936.4]
  wire  _T_12862; // @[Mux.scala 46:19:@10937.4]
  wire [7:0] _T_12863; // @[Mux.scala 46:16:@10938.4]
  wire  _T_12864; // @[Mux.scala 46:19:@10939.4]
  wire [7:0] _T_12865; // @[Mux.scala 46:16:@10940.4]
  wire  _T_12866; // @[Mux.scala 46:19:@10941.4]
  wire [7:0] _T_12867; // @[Mux.scala 46:16:@10942.4]
  wire  _T_12868; // @[Mux.scala 46:19:@10943.4]
  wire [7:0] _T_12869; // @[Mux.scala 46:16:@10944.4]
  wire  _T_12870; // @[Mux.scala 46:19:@10945.4]
  wire [7:0] _T_12871; // @[Mux.scala 46:16:@10946.4]
  wire  _T_12872; // @[Mux.scala 46:19:@10947.4]
  wire [7:0] _T_12873; // @[Mux.scala 46:16:@10948.4]
  wire  _T_12874; // @[Mux.scala 46:19:@10949.4]
  wire [7:0] _T_12875; // @[Mux.scala 46:16:@10950.4]
  wire  _T_12876; // @[Mux.scala 46:19:@10951.4]
  wire [7:0] _T_12877; // @[Mux.scala 46:16:@10952.4]
  wire  _T_12878; // @[Mux.scala 46:19:@10953.4]
  wire [7:0] _T_12879; // @[Mux.scala 46:16:@10954.4]
  wire  _T_12880; // @[Mux.scala 46:19:@10955.4]
  wire [7:0] _T_12881; // @[Mux.scala 46:16:@10956.4]
  wire  _T_12882; // @[Mux.scala 46:19:@10957.4]
  wire [7:0] _T_12883; // @[Mux.scala 46:16:@10958.4]
  wire  _T_12884; // @[Mux.scala 46:19:@10959.4]
  wire [7:0] _T_12885; // @[Mux.scala 46:16:@10960.4]
  wire  _T_12886; // @[Mux.scala 46:19:@10961.4]
  wire [7:0] _T_12887; // @[Mux.scala 46:16:@10962.4]
  wire  _T_12888; // @[Mux.scala 46:19:@10963.4]
  wire [7:0] _T_12889; // @[Mux.scala 46:16:@10964.4]
  wire  _T_12890; // @[Mux.scala 46:19:@10965.4]
  wire [7:0] _T_12891; // @[Mux.scala 46:16:@10966.4]
  wire  _T_12892; // @[Mux.scala 46:19:@10967.4]
  wire [7:0] _T_12893; // @[Mux.scala 46:16:@10968.4]
  wire  _T_12894; // @[Mux.scala 46:19:@10969.4]
  wire [7:0] _T_12895; // @[Mux.scala 46:16:@10970.4]
  wire  _T_12896; // @[Mux.scala 46:19:@10971.4]
  wire [7:0] _T_12897; // @[Mux.scala 46:16:@10972.4]
  wire  _T_12898; // @[Mux.scala 46:19:@10973.4]
  wire [7:0] _T_12899; // @[Mux.scala 46:16:@10974.4]
  wire  _T_12900; // @[Mux.scala 46:19:@10975.4]
  wire [7:0] _T_12901; // @[Mux.scala 46:16:@10976.4]
  wire  _T_12902; // @[Mux.scala 46:19:@10977.4]
  wire [7:0] _T_12903; // @[Mux.scala 46:16:@10978.4]
  wire  _T_12904; // @[Mux.scala 46:19:@10979.4]
  wire [7:0] _T_12905; // @[Mux.scala 46:16:@10980.4]
  wire  _T_12906; // @[Mux.scala 46:19:@10981.4]
  wire [7:0] _T_12907; // @[Mux.scala 46:16:@10982.4]
  wire  _T_12908; // @[Mux.scala 46:19:@10983.4]
  wire [7:0] _T_12909; // @[Mux.scala 46:16:@10984.4]
  wire  _T_12952; // @[Mux.scala 46:19:@10986.4]
  wire [7:0] _T_12953; // @[Mux.scala 46:16:@10987.4]
  wire  _T_12954; // @[Mux.scala 46:19:@10988.4]
  wire [7:0] _T_12955; // @[Mux.scala 46:16:@10989.4]
  wire  _T_12956; // @[Mux.scala 46:19:@10990.4]
  wire [7:0] _T_12957; // @[Mux.scala 46:16:@10991.4]
  wire  _T_12958; // @[Mux.scala 46:19:@10992.4]
  wire [7:0] _T_12959; // @[Mux.scala 46:16:@10993.4]
  wire  _T_12960; // @[Mux.scala 46:19:@10994.4]
  wire [7:0] _T_12961; // @[Mux.scala 46:16:@10995.4]
  wire  _T_12962; // @[Mux.scala 46:19:@10996.4]
  wire [7:0] _T_12963; // @[Mux.scala 46:16:@10997.4]
  wire  _T_12964; // @[Mux.scala 46:19:@10998.4]
  wire [7:0] _T_12965; // @[Mux.scala 46:16:@10999.4]
  wire  _T_12966; // @[Mux.scala 46:19:@11000.4]
  wire [7:0] _T_12967; // @[Mux.scala 46:16:@11001.4]
  wire  _T_12968; // @[Mux.scala 46:19:@11002.4]
  wire [7:0] _T_12969; // @[Mux.scala 46:16:@11003.4]
  wire  _T_12970; // @[Mux.scala 46:19:@11004.4]
  wire [7:0] _T_12971; // @[Mux.scala 46:16:@11005.4]
  wire  _T_12972; // @[Mux.scala 46:19:@11006.4]
  wire [7:0] _T_12973; // @[Mux.scala 46:16:@11007.4]
  wire  _T_12974; // @[Mux.scala 46:19:@11008.4]
  wire [7:0] _T_12975; // @[Mux.scala 46:16:@11009.4]
  wire  _T_12976; // @[Mux.scala 46:19:@11010.4]
  wire [7:0] _T_12977; // @[Mux.scala 46:16:@11011.4]
  wire  _T_12978; // @[Mux.scala 46:19:@11012.4]
  wire [7:0] _T_12979; // @[Mux.scala 46:16:@11013.4]
  wire  _T_12980; // @[Mux.scala 46:19:@11014.4]
  wire [7:0] _T_12981; // @[Mux.scala 46:16:@11015.4]
  wire  _T_12982; // @[Mux.scala 46:19:@11016.4]
  wire [7:0] _T_12983; // @[Mux.scala 46:16:@11017.4]
  wire  _T_12984; // @[Mux.scala 46:19:@11018.4]
  wire [7:0] _T_12985; // @[Mux.scala 46:16:@11019.4]
  wire  _T_12986; // @[Mux.scala 46:19:@11020.4]
  wire [7:0] _T_12987; // @[Mux.scala 46:16:@11021.4]
  wire  _T_12988; // @[Mux.scala 46:19:@11022.4]
  wire [7:0] _T_12989; // @[Mux.scala 46:16:@11023.4]
  wire  _T_12990; // @[Mux.scala 46:19:@11024.4]
  wire [7:0] _T_12991; // @[Mux.scala 46:16:@11025.4]
  wire  _T_12992; // @[Mux.scala 46:19:@11026.4]
  wire [7:0] _T_12993; // @[Mux.scala 46:16:@11027.4]
  wire  _T_12994; // @[Mux.scala 46:19:@11028.4]
  wire [7:0] _T_12995; // @[Mux.scala 46:16:@11029.4]
  wire  _T_12996; // @[Mux.scala 46:19:@11030.4]
  wire [7:0] _T_12997; // @[Mux.scala 46:16:@11031.4]
  wire  _T_12998; // @[Mux.scala 46:19:@11032.4]
  wire [7:0] _T_12999; // @[Mux.scala 46:16:@11033.4]
  wire  _T_13000; // @[Mux.scala 46:19:@11034.4]
  wire [7:0] _T_13001; // @[Mux.scala 46:16:@11035.4]
  wire  _T_13002; // @[Mux.scala 46:19:@11036.4]
  wire [7:0] _T_13003; // @[Mux.scala 46:16:@11037.4]
  wire  _T_13004; // @[Mux.scala 46:19:@11038.4]
  wire [7:0] _T_13005; // @[Mux.scala 46:16:@11039.4]
  wire  _T_13006; // @[Mux.scala 46:19:@11040.4]
  wire [7:0] _T_13007; // @[Mux.scala 46:16:@11041.4]
  wire  _T_13008; // @[Mux.scala 46:19:@11042.4]
  wire [7:0] _T_13009; // @[Mux.scala 46:16:@11043.4]
  wire  _T_13010; // @[Mux.scala 46:19:@11044.4]
  wire [7:0] _T_13011; // @[Mux.scala 46:16:@11045.4]
  wire  _T_13012; // @[Mux.scala 46:19:@11046.4]
  wire [7:0] _T_13013; // @[Mux.scala 46:16:@11047.4]
  wire  _T_13014; // @[Mux.scala 46:19:@11048.4]
  wire [7:0] _T_13015; // @[Mux.scala 46:16:@11049.4]
  wire  _T_13016; // @[Mux.scala 46:19:@11050.4]
  wire [7:0] _T_13017; // @[Mux.scala 46:16:@11051.4]
  wire  _T_13018; // @[Mux.scala 46:19:@11052.4]
  wire [7:0] _T_13019; // @[Mux.scala 46:16:@11053.4]
  wire  _T_13020; // @[Mux.scala 46:19:@11054.4]
  wire [7:0] _T_13021; // @[Mux.scala 46:16:@11055.4]
  wire  _T_13022; // @[Mux.scala 46:19:@11056.4]
  wire [7:0] _T_13023; // @[Mux.scala 46:16:@11057.4]
  wire  _T_13024; // @[Mux.scala 46:19:@11058.4]
  wire [7:0] _T_13025; // @[Mux.scala 46:16:@11059.4]
  wire  _T_13026; // @[Mux.scala 46:19:@11060.4]
  wire [7:0] _T_13027; // @[Mux.scala 46:16:@11061.4]
  wire  _T_13028; // @[Mux.scala 46:19:@11062.4]
  wire [7:0] _T_13029; // @[Mux.scala 46:16:@11063.4]
  wire  _T_13030; // @[Mux.scala 46:19:@11064.4]
  wire [7:0] _T_13031; // @[Mux.scala 46:16:@11065.4]
  wire  _T_13032; // @[Mux.scala 46:19:@11066.4]
  wire [7:0] _T_13033; // @[Mux.scala 46:16:@11067.4]
  wire  _T_13077; // @[Mux.scala 46:19:@11069.4]
  wire [7:0] _T_13078; // @[Mux.scala 46:16:@11070.4]
  wire  _T_13079; // @[Mux.scala 46:19:@11071.4]
  wire [7:0] _T_13080; // @[Mux.scala 46:16:@11072.4]
  wire  _T_13081; // @[Mux.scala 46:19:@11073.4]
  wire [7:0] _T_13082; // @[Mux.scala 46:16:@11074.4]
  wire  _T_13083; // @[Mux.scala 46:19:@11075.4]
  wire [7:0] _T_13084; // @[Mux.scala 46:16:@11076.4]
  wire  _T_13085; // @[Mux.scala 46:19:@11077.4]
  wire [7:0] _T_13086; // @[Mux.scala 46:16:@11078.4]
  wire  _T_13087; // @[Mux.scala 46:19:@11079.4]
  wire [7:0] _T_13088; // @[Mux.scala 46:16:@11080.4]
  wire  _T_13089; // @[Mux.scala 46:19:@11081.4]
  wire [7:0] _T_13090; // @[Mux.scala 46:16:@11082.4]
  wire  _T_13091; // @[Mux.scala 46:19:@11083.4]
  wire [7:0] _T_13092; // @[Mux.scala 46:16:@11084.4]
  wire  _T_13093; // @[Mux.scala 46:19:@11085.4]
  wire [7:0] _T_13094; // @[Mux.scala 46:16:@11086.4]
  wire  _T_13095; // @[Mux.scala 46:19:@11087.4]
  wire [7:0] _T_13096; // @[Mux.scala 46:16:@11088.4]
  wire  _T_13097; // @[Mux.scala 46:19:@11089.4]
  wire [7:0] _T_13098; // @[Mux.scala 46:16:@11090.4]
  wire  _T_13099; // @[Mux.scala 46:19:@11091.4]
  wire [7:0] _T_13100; // @[Mux.scala 46:16:@11092.4]
  wire  _T_13101; // @[Mux.scala 46:19:@11093.4]
  wire [7:0] _T_13102; // @[Mux.scala 46:16:@11094.4]
  wire  _T_13103; // @[Mux.scala 46:19:@11095.4]
  wire [7:0] _T_13104; // @[Mux.scala 46:16:@11096.4]
  wire  _T_13105; // @[Mux.scala 46:19:@11097.4]
  wire [7:0] _T_13106; // @[Mux.scala 46:16:@11098.4]
  wire  _T_13107; // @[Mux.scala 46:19:@11099.4]
  wire [7:0] _T_13108; // @[Mux.scala 46:16:@11100.4]
  wire  _T_13109; // @[Mux.scala 46:19:@11101.4]
  wire [7:0] _T_13110; // @[Mux.scala 46:16:@11102.4]
  wire  _T_13111; // @[Mux.scala 46:19:@11103.4]
  wire [7:0] _T_13112; // @[Mux.scala 46:16:@11104.4]
  wire  _T_13113; // @[Mux.scala 46:19:@11105.4]
  wire [7:0] _T_13114; // @[Mux.scala 46:16:@11106.4]
  wire  _T_13115; // @[Mux.scala 46:19:@11107.4]
  wire [7:0] _T_13116; // @[Mux.scala 46:16:@11108.4]
  wire  _T_13117; // @[Mux.scala 46:19:@11109.4]
  wire [7:0] _T_13118; // @[Mux.scala 46:16:@11110.4]
  wire  _T_13119; // @[Mux.scala 46:19:@11111.4]
  wire [7:0] _T_13120; // @[Mux.scala 46:16:@11112.4]
  wire  _T_13121; // @[Mux.scala 46:19:@11113.4]
  wire [7:0] _T_13122; // @[Mux.scala 46:16:@11114.4]
  wire  _T_13123; // @[Mux.scala 46:19:@11115.4]
  wire [7:0] _T_13124; // @[Mux.scala 46:16:@11116.4]
  wire  _T_13125; // @[Mux.scala 46:19:@11117.4]
  wire [7:0] _T_13126; // @[Mux.scala 46:16:@11118.4]
  wire  _T_13127; // @[Mux.scala 46:19:@11119.4]
  wire [7:0] _T_13128; // @[Mux.scala 46:16:@11120.4]
  wire  _T_13129; // @[Mux.scala 46:19:@11121.4]
  wire [7:0] _T_13130; // @[Mux.scala 46:16:@11122.4]
  wire  _T_13131; // @[Mux.scala 46:19:@11123.4]
  wire [7:0] _T_13132; // @[Mux.scala 46:16:@11124.4]
  wire  _T_13133; // @[Mux.scala 46:19:@11125.4]
  wire [7:0] _T_13134; // @[Mux.scala 46:16:@11126.4]
  wire  _T_13135; // @[Mux.scala 46:19:@11127.4]
  wire [7:0] _T_13136; // @[Mux.scala 46:16:@11128.4]
  wire  _T_13137; // @[Mux.scala 46:19:@11129.4]
  wire [7:0] _T_13138; // @[Mux.scala 46:16:@11130.4]
  wire  _T_13139; // @[Mux.scala 46:19:@11131.4]
  wire [7:0] _T_13140; // @[Mux.scala 46:16:@11132.4]
  wire  _T_13141; // @[Mux.scala 46:19:@11133.4]
  wire [7:0] _T_13142; // @[Mux.scala 46:16:@11134.4]
  wire  _T_13143; // @[Mux.scala 46:19:@11135.4]
  wire [7:0] _T_13144; // @[Mux.scala 46:16:@11136.4]
  wire  _T_13145; // @[Mux.scala 46:19:@11137.4]
  wire [7:0] _T_13146; // @[Mux.scala 46:16:@11138.4]
  wire  _T_13147; // @[Mux.scala 46:19:@11139.4]
  wire [7:0] _T_13148; // @[Mux.scala 46:16:@11140.4]
  wire  _T_13149; // @[Mux.scala 46:19:@11141.4]
  wire [7:0] _T_13150; // @[Mux.scala 46:16:@11142.4]
  wire  _T_13151; // @[Mux.scala 46:19:@11143.4]
  wire [7:0] _T_13152; // @[Mux.scala 46:16:@11144.4]
  wire  _T_13153; // @[Mux.scala 46:19:@11145.4]
  wire [7:0] _T_13154; // @[Mux.scala 46:16:@11146.4]
  wire  _T_13155; // @[Mux.scala 46:19:@11147.4]
  wire [7:0] _T_13156; // @[Mux.scala 46:16:@11148.4]
  wire  _T_13157; // @[Mux.scala 46:19:@11149.4]
  wire [7:0] _T_13158; // @[Mux.scala 46:16:@11150.4]
  wire  _T_13159; // @[Mux.scala 46:19:@11151.4]
  wire [7:0] _T_13160; // @[Mux.scala 46:16:@11152.4]
  wire  _T_13205; // @[Mux.scala 46:19:@11154.4]
  wire [7:0] _T_13206; // @[Mux.scala 46:16:@11155.4]
  wire  _T_13207; // @[Mux.scala 46:19:@11156.4]
  wire [7:0] _T_13208; // @[Mux.scala 46:16:@11157.4]
  wire  _T_13209; // @[Mux.scala 46:19:@11158.4]
  wire [7:0] _T_13210; // @[Mux.scala 46:16:@11159.4]
  wire  _T_13211; // @[Mux.scala 46:19:@11160.4]
  wire [7:0] _T_13212; // @[Mux.scala 46:16:@11161.4]
  wire  _T_13213; // @[Mux.scala 46:19:@11162.4]
  wire [7:0] _T_13214; // @[Mux.scala 46:16:@11163.4]
  wire  _T_13215; // @[Mux.scala 46:19:@11164.4]
  wire [7:0] _T_13216; // @[Mux.scala 46:16:@11165.4]
  wire  _T_13217; // @[Mux.scala 46:19:@11166.4]
  wire [7:0] _T_13218; // @[Mux.scala 46:16:@11167.4]
  wire  _T_13219; // @[Mux.scala 46:19:@11168.4]
  wire [7:0] _T_13220; // @[Mux.scala 46:16:@11169.4]
  wire  _T_13221; // @[Mux.scala 46:19:@11170.4]
  wire [7:0] _T_13222; // @[Mux.scala 46:16:@11171.4]
  wire  _T_13223; // @[Mux.scala 46:19:@11172.4]
  wire [7:0] _T_13224; // @[Mux.scala 46:16:@11173.4]
  wire  _T_13225; // @[Mux.scala 46:19:@11174.4]
  wire [7:0] _T_13226; // @[Mux.scala 46:16:@11175.4]
  wire  _T_13227; // @[Mux.scala 46:19:@11176.4]
  wire [7:0] _T_13228; // @[Mux.scala 46:16:@11177.4]
  wire  _T_13229; // @[Mux.scala 46:19:@11178.4]
  wire [7:0] _T_13230; // @[Mux.scala 46:16:@11179.4]
  wire  _T_13231; // @[Mux.scala 46:19:@11180.4]
  wire [7:0] _T_13232; // @[Mux.scala 46:16:@11181.4]
  wire  _T_13233; // @[Mux.scala 46:19:@11182.4]
  wire [7:0] _T_13234; // @[Mux.scala 46:16:@11183.4]
  wire  _T_13235; // @[Mux.scala 46:19:@11184.4]
  wire [7:0] _T_13236; // @[Mux.scala 46:16:@11185.4]
  wire  _T_13237; // @[Mux.scala 46:19:@11186.4]
  wire [7:0] _T_13238; // @[Mux.scala 46:16:@11187.4]
  wire  _T_13239; // @[Mux.scala 46:19:@11188.4]
  wire [7:0] _T_13240; // @[Mux.scala 46:16:@11189.4]
  wire  _T_13241; // @[Mux.scala 46:19:@11190.4]
  wire [7:0] _T_13242; // @[Mux.scala 46:16:@11191.4]
  wire  _T_13243; // @[Mux.scala 46:19:@11192.4]
  wire [7:0] _T_13244; // @[Mux.scala 46:16:@11193.4]
  wire  _T_13245; // @[Mux.scala 46:19:@11194.4]
  wire [7:0] _T_13246; // @[Mux.scala 46:16:@11195.4]
  wire  _T_13247; // @[Mux.scala 46:19:@11196.4]
  wire [7:0] _T_13248; // @[Mux.scala 46:16:@11197.4]
  wire  _T_13249; // @[Mux.scala 46:19:@11198.4]
  wire [7:0] _T_13250; // @[Mux.scala 46:16:@11199.4]
  wire  _T_13251; // @[Mux.scala 46:19:@11200.4]
  wire [7:0] _T_13252; // @[Mux.scala 46:16:@11201.4]
  wire  _T_13253; // @[Mux.scala 46:19:@11202.4]
  wire [7:0] _T_13254; // @[Mux.scala 46:16:@11203.4]
  wire  _T_13255; // @[Mux.scala 46:19:@11204.4]
  wire [7:0] _T_13256; // @[Mux.scala 46:16:@11205.4]
  wire  _T_13257; // @[Mux.scala 46:19:@11206.4]
  wire [7:0] _T_13258; // @[Mux.scala 46:16:@11207.4]
  wire  _T_13259; // @[Mux.scala 46:19:@11208.4]
  wire [7:0] _T_13260; // @[Mux.scala 46:16:@11209.4]
  wire  _T_13261; // @[Mux.scala 46:19:@11210.4]
  wire [7:0] _T_13262; // @[Mux.scala 46:16:@11211.4]
  wire  _T_13263; // @[Mux.scala 46:19:@11212.4]
  wire [7:0] _T_13264; // @[Mux.scala 46:16:@11213.4]
  wire  _T_13265; // @[Mux.scala 46:19:@11214.4]
  wire [7:0] _T_13266; // @[Mux.scala 46:16:@11215.4]
  wire  _T_13267; // @[Mux.scala 46:19:@11216.4]
  wire [7:0] _T_13268; // @[Mux.scala 46:16:@11217.4]
  wire  _T_13269; // @[Mux.scala 46:19:@11218.4]
  wire [7:0] _T_13270; // @[Mux.scala 46:16:@11219.4]
  wire  _T_13271; // @[Mux.scala 46:19:@11220.4]
  wire [7:0] _T_13272; // @[Mux.scala 46:16:@11221.4]
  wire  _T_13273; // @[Mux.scala 46:19:@11222.4]
  wire [7:0] _T_13274; // @[Mux.scala 46:16:@11223.4]
  wire  _T_13275; // @[Mux.scala 46:19:@11224.4]
  wire [7:0] _T_13276; // @[Mux.scala 46:16:@11225.4]
  wire  _T_13277; // @[Mux.scala 46:19:@11226.4]
  wire [7:0] _T_13278; // @[Mux.scala 46:16:@11227.4]
  wire  _T_13279; // @[Mux.scala 46:19:@11228.4]
  wire [7:0] _T_13280; // @[Mux.scala 46:16:@11229.4]
  wire  _T_13281; // @[Mux.scala 46:19:@11230.4]
  wire [7:0] _T_13282; // @[Mux.scala 46:16:@11231.4]
  wire  _T_13283; // @[Mux.scala 46:19:@11232.4]
  wire [7:0] _T_13284; // @[Mux.scala 46:16:@11233.4]
  wire  _T_13285; // @[Mux.scala 46:19:@11234.4]
  wire [7:0] _T_13286; // @[Mux.scala 46:16:@11235.4]
  wire  _T_13287; // @[Mux.scala 46:19:@11236.4]
  wire [7:0] _T_13288; // @[Mux.scala 46:16:@11237.4]
  wire  _T_13289; // @[Mux.scala 46:19:@11238.4]
  wire [7:0] _T_13290; // @[Mux.scala 46:16:@11239.4]
  wire  _T_13336; // @[Mux.scala 46:19:@11241.4]
  wire [7:0] _T_13337; // @[Mux.scala 46:16:@11242.4]
  wire  _T_13338; // @[Mux.scala 46:19:@11243.4]
  wire [7:0] _T_13339; // @[Mux.scala 46:16:@11244.4]
  wire  _T_13340; // @[Mux.scala 46:19:@11245.4]
  wire [7:0] _T_13341; // @[Mux.scala 46:16:@11246.4]
  wire  _T_13342; // @[Mux.scala 46:19:@11247.4]
  wire [7:0] _T_13343; // @[Mux.scala 46:16:@11248.4]
  wire  _T_13344; // @[Mux.scala 46:19:@11249.4]
  wire [7:0] _T_13345; // @[Mux.scala 46:16:@11250.4]
  wire  _T_13346; // @[Mux.scala 46:19:@11251.4]
  wire [7:0] _T_13347; // @[Mux.scala 46:16:@11252.4]
  wire  _T_13348; // @[Mux.scala 46:19:@11253.4]
  wire [7:0] _T_13349; // @[Mux.scala 46:16:@11254.4]
  wire  _T_13350; // @[Mux.scala 46:19:@11255.4]
  wire [7:0] _T_13351; // @[Mux.scala 46:16:@11256.4]
  wire  _T_13352; // @[Mux.scala 46:19:@11257.4]
  wire [7:0] _T_13353; // @[Mux.scala 46:16:@11258.4]
  wire  _T_13354; // @[Mux.scala 46:19:@11259.4]
  wire [7:0] _T_13355; // @[Mux.scala 46:16:@11260.4]
  wire  _T_13356; // @[Mux.scala 46:19:@11261.4]
  wire [7:0] _T_13357; // @[Mux.scala 46:16:@11262.4]
  wire  _T_13358; // @[Mux.scala 46:19:@11263.4]
  wire [7:0] _T_13359; // @[Mux.scala 46:16:@11264.4]
  wire  _T_13360; // @[Mux.scala 46:19:@11265.4]
  wire [7:0] _T_13361; // @[Mux.scala 46:16:@11266.4]
  wire  _T_13362; // @[Mux.scala 46:19:@11267.4]
  wire [7:0] _T_13363; // @[Mux.scala 46:16:@11268.4]
  wire  _T_13364; // @[Mux.scala 46:19:@11269.4]
  wire [7:0] _T_13365; // @[Mux.scala 46:16:@11270.4]
  wire  _T_13366; // @[Mux.scala 46:19:@11271.4]
  wire [7:0] _T_13367; // @[Mux.scala 46:16:@11272.4]
  wire  _T_13368; // @[Mux.scala 46:19:@11273.4]
  wire [7:0] _T_13369; // @[Mux.scala 46:16:@11274.4]
  wire  _T_13370; // @[Mux.scala 46:19:@11275.4]
  wire [7:0] _T_13371; // @[Mux.scala 46:16:@11276.4]
  wire  _T_13372; // @[Mux.scala 46:19:@11277.4]
  wire [7:0] _T_13373; // @[Mux.scala 46:16:@11278.4]
  wire  _T_13374; // @[Mux.scala 46:19:@11279.4]
  wire [7:0] _T_13375; // @[Mux.scala 46:16:@11280.4]
  wire  _T_13376; // @[Mux.scala 46:19:@11281.4]
  wire [7:0] _T_13377; // @[Mux.scala 46:16:@11282.4]
  wire  _T_13378; // @[Mux.scala 46:19:@11283.4]
  wire [7:0] _T_13379; // @[Mux.scala 46:16:@11284.4]
  wire  _T_13380; // @[Mux.scala 46:19:@11285.4]
  wire [7:0] _T_13381; // @[Mux.scala 46:16:@11286.4]
  wire  _T_13382; // @[Mux.scala 46:19:@11287.4]
  wire [7:0] _T_13383; // @[Mux.scala 46:16:@11288.4]
  wire  _T_13384; // @[Mux.scala 46:19:@11289.4]
  wire [7:0] _T_13385; // @[Mux.scala 46:16:@11290.4]
  wire  _T_13386; // @[Mux.scala 46:19:@11291.4]
  wire [7:0] _T_13387; // @[Mux.scala 46:16:@11292.4]
  wire  _T_13388; // @[Mux.scala 46:19:@11293.4]
  wire [7:0] _T_13389; // @[Mux.scala 46:16:@11294.4]
  wire  _T_13390; // @[Mux.scala 46:19:@11295.4]
  wire [7:0] _T_13391; // @[Mux.scala 46:16:@11296.4]
  wire  _T_13392; // @[Mux.scala 46:19:@11297.4]
  wire [7:0] _T_13393; // @[Mux.scala 46:16:@11298.4]
  wire  _T_13394; // @[Mux.scala 46:19:@11299.4]
  wire [7:0] _T_13395; // @[Mux.scala 46:16:@11300.4]
  wire  _T_13396; // @[Mux.scala 46:19:@11301.4]
  wire [7:0] _T_13397; // @[Mux.scala 46:16:@11302.4]
  wire  _T_13398; // @[Mux.scala 46:19:@11303.4]
  wire [7:0] _T_13399; // @[Mux.scala 46:16:@11304.4]
  wire  _T_13400; // @[Mux.scala 46:19:@11305.4]
  wire [7:0] _T_13401; // @[Mux.scala 46:16:@11306.4]
  wire  _T_13402; // @[Mux.scala 46:19:@11307.4]
  wire [7:0] _T_13403; // @[Mux.scala 46:16:@11308.4]
  wire  _T_13404; // @[Mux.scala 46:19:@11309.4]
  wire [7:0] _T_13405; // @[Mux.scala 46:16:@11310.4]
  wire  _T_13406; // @[Mux.scala 46:19:@11311.4]
  wire [7:0] _T_13407; // @[Mux.scala 46:16:@11312.4]
  wire  _T_13408; // @[Mux.scala 46:19:@11313.4]
  wire [7:0] _T_13409; // @[Mux.scala 46:16:@11314.4]
  wire  _T_13410; // @[Mux.scala 46:19:@11315.4]
  wire [7:0] _T_13411; // @[Mux.scala 46:16:@11316.4]
  wire  _T_13412; // @[Mux.scala 46:19:@11317.4]
  wire [7:0] _T_13413; // @[Mux.scala 46:16:@11318.4]
  wire  _T_13414; // @[Mux.scala 46:19:@11319.4]
  wire [7:0] _T_13415; // @[Mux.scala 46:16:@11320.4]
  wire  _T_13416; // @[Mux.scala 46:19:@11321.4]
  wire [7:0] _T_13417; // @[Mux.scala 46:16:@11322.4]
  wire  _T_13418; // @[Mux.scala 46:19:@11323.4]
  wire [7:0] _T_13419; // @[Mux.scala 46:16:@11324.4]
  wire  _T_13420; // @[Mux.scala 46:19:@11325.4]
  wire [7:0] _T_13421; // @[Mux.scala 46:16:@11326.4]
  wire  _T_13422; // @[Mux.scala 46:19:@11327.4]
  wire [7:0] _T_13423; // @[Mux.scala 46:16:@11328.4]
  wire  _T_13470; // @[Mux.scala 46:19:@11330.4]
  wire [7:0] _T_13471; // @[Mux.scala 46:16:@11331.4]
  wire  _T_13472; // @[Mux.scala 46:19:@11332.4]
  wire [7:0] _T_13473; // @[Mux.scala 46:16:@11333.4]
  wire  _T_13474; // @[Mux.scala 46:19:@11334.4]
  wire [7:0] _T_13475; // @[Mux.scala 46:16:@11335.4]
  wire  _T_13476; // @[Mux.scala 46:19:@11336.4]
  wire [7:0] _T_13477; // @[Mux.scala 46:16:@11337.4]
  wire  _T_13478; // @[Mux.scala 46:19:@11338.4]
  wire [7:0] _T_13479; // @[Mux.scala 46:16:@11339.4]
  wire  _T_13480; // @[Mux.scala 46:19:@11340.4]
  wire [7:0] _T_13481; // @[Mux.scala 46:16:@11341.4]
  wire  _T_13482; // @[Mux.scala 46:19:@11342.4]
  wire [7:0] _T_13483; // @[Mux.scala 46:16:@11343.4]
  wire  _T_13484; // @[Mux.scala 46:19:@11344.4]
  wire [7:0] _T_13485; // @[Mux.scala 46:16:@11345.4]
  wire  _T_13486; // @[Mux.scala 46:19:@11346.4]
  wire [7:0] _T_13487; // @[Mux.scala 46:16:@11347.4]
  wire  _T_13488; // @[Mux.scala 46:19:@11348.4]
  wire [7:0] _T_13489; // @[Mux.scala 46:16:@11349.4]
  wire  _T_13490; // @[Mux.scala 46:19:@11350.4]
  wire [7:0] _T_13491; // @[Mux.scala 46:16:@11351.4]
  wire  _T_13492; // @[Mux.scala 46:19:@11352.4]
  wire [7:0] _T_13493; // @[Mux.scala 46:16:@11353.4]
  wire  _T_13494; // @[Mux.scala 46:19:@11354.4]
  wire [7:0] _T_13495; // @[Mux.scala 46:16:@11355.4]
  wire  _T_13496; // @[Mux.scala 46:19:@11356.4]
  wire [7:0] _T_13497; // @[Mux.scala 46:16:@11357.4]
  wire  _T_13498; // @[Mux.scala 46:19:@11358.4]
  wire [7:0] _T_13499; // @[Mux.scala 46:16:@11359.4]
  wire  _T_13500; // @[Mux.scala 46:19:@11360.4]
  wire [7:0] _T_13501; // @[Mux.scala 46:16:@11361.4]
  wire  _T_13502; // @[Mux.scala 46:19:@11362.4]
  wire [7:0] _T_13503; // @[Mux.scala 46:16:@11363.4]
  wire  _T_13504; // @[Mux.scala 46:19:@11364.4]
  wire [7:0] _T_13505; // @[Mux.scala 46:16:@11365.4]
  wire  _T_13506; // @[Mux.scala 46:19:@11366.4]
  wire [7:0] _T_13507; // @[Mux.scala 46:16:@11367.4]
  wire  _T_13508; // @[Mux.scala 46:19:@11368.4]
  wire [7:0] _T_13509; // @[Mux.scala 46:16:@11369.4]
  wire  _T_13510; // @[Mux.scala 46:19:@11370.4]
  wire [7:0] _T_13511; // @[Mux.scala 46:16:@11371.4]
  wire  _T_13512; // @[Mux.scala 46:19:@11372.4]
  wire [7:0] _T_13513; // @[Mux.scala 46:16:@11373.4]
  wire  _T_13514; // @[Mux.scala 46:19:@11374.4]
  wire [7:0] _T_13515; // @[Mux.scala 46:16:@11375.4]
  wire  _T_13516; // @[Mux.scala 46:19:@11376.4]
  wire [7:0] _T_13517; // @[Mux.scala 46:16:@11377.4]
  wire  _T_13518; // @[Mux.scala 46:19:@11378.4]
  wire [7:0] _T_13519; // @[Mux.scala 46:16:@11379.4]
  wire  _T_13520; // @[Mux.scala 46:19:@11380.4]
  wire [7:0] _T_13521; // @[Mux.scala 46:16:@11381.4]
  wire  _T_13522; // @[Mux.scala 46:19:@11382.4]
  wire [7:0] _T_13523; // @[Mux.scala 46:16:@11383.4]
  wire  _T_13524; // @[Mux.scala 46:19:@11384.4]
  wire [7:0] _T_13525; // @[Mux.scala 46:16:@11385.4]
  wire  _T_13526; // @[Mux.scala 46:19:@11386.4]
  wire [7:0] _T_13527; // @[Mux.scala 46:16:@11387.4]
  wire  _T_13528; // @[Mux.scala 46:19:@11388.4]
  wire [7:0] _T_13529; // @[Mux.scala 46:16:@11389.4]
  wire  _T_13530; // @[Mux.scala 46:19:@11390.4]
  wire [7:0] _T_13531; // @[Mux.scala 46:16:@11391.4]
  wire  _T_13532; // @[Mux.scala 46:19:@11392.4]
  wire [7:0] _T_13533; // @[Mux.scala 46:16:@11393.4]
  wire  _T_13534; // @[Mux.scala 46:19:@11394.4]
  wire [7:0] _T_13535; // @[Mux.scala 46:16:@11395.4]
  wire  _T_13536; // @[Mux.scala 46:19:@11396.4]
  wire [7:0] _T_13537; // @[Mux.scala 46:16:@11397.4]
  wire  _T_13538; // @[Mux.scala 46:19:@11398.4]
  wire [7:0] _T_13539; // @[Mux.scala 46:16:@11399.4]
  wire  _T_13540; // @[Mux.scala 46:19:@11400.4]
  wire [7:0] _T_13541; // @[Mux.scala 46:16:@11401.4]
  wire  _T_13542; // @[Mux.scala 46:19:@11402.4]
  wire [7:0] _T_13543; // @[Mux.scala 46:16:@11403.4]
  wire  _T_13544; // @[Mux.scala 46:19:@11404.4]
  wire [7:0] _T_13545; // @[Mux.scala 46:16:@11405.4]
  wire  _T_13546; // @[Mux.scala 46:19:@11406.4]
  wire [7:0] _T_13547; // @[Mux.scala 46:16:@11407.4]
  wire  _T_13548; // @[Mux.scala 46:19:@11408.4]
  wire [7:0] _T_13549; // @[Mux.scala 46:16:@11409.4]
  wire  _T_13550; // @[Mux.scala 46:19:@11410.4]
  wire [7:0] _T_13551; // @[Mux.scala 46:16:@11411.4]
  wire  _T_13552; // @[Mux.scala 46:19:@11412.4]
  wire [7:0] _T_13553; // @[Mux.scala 46:16:@11413.4]
  wire  _T_13554; // @[Mux.scala 46:19:@11414.4]
  wire [7:0] _T_13555; // @[Mux.scala 46:16:@11415.4]
  wire  _T_13556; // @[Mux.scala 46:19:@11416.4]
  wire [7:0] _T_13557; // @[Mux.scala 46:16:@11417.4]
  wire  _T_13558; // @[Mux.scala 46:19:@11418.4]
  wire [7:0] _T_13559; // @[Mux.scala 46:16:@11419.4]
  wire  _T_13607; // @[Mux.scala 46:19:@11421.4]
  wire [7:0] _T_13608; // @[Mux.scala 46:16:@11422.4]
  wire  _T_13609; // @[Mux.scala 46:19:@11423.4]
  wire [7:0] _T_13610; // @[Mux.scala 46:16:@11424.4]
  wire  _T_13611; // @[Mux.scala 46:19:@11425.4]
  wire [7:0] _T_13612; // @[Mux.scala 46:16:@11426.4]
  wire  _T_13613; // @[Mux.scala 46:19:@11427.4]
  wire [7:0] _T_13614; // @[Mux.scala 46:16:@11428.4]
  wire  _T_13615; // @[Mux.scala 46:19:@11429.4]
  wire [7:0] _T_13616; // @[Mux.scala 46:16:@11430.4]
  wire  _T_13617; // @[Mux.scala 46:19:@11431.4]
  wire [7:0] _T_13618; // @[Mux.scala 46:16:@11432.4]
  wire  _T_13619; // @[Mux.scala 46:19:@11433.4]
  wire [7:0] _T_13620; // @[Mux.scala 46:16:@11434.4]
  wire  _T_13621; // @[Mux.scala 46:19:@11435.4]
  wire [7:0] _T_13622; // @[Mux.scala 46:16:@11436.4]
  wire  _T_13623; // @[Mux.scala 46:19:@11437.4]
  wire [7:0] _T_13624; // @[Mux.scala 46:16:@11438.4]
  wire  _T_13625; // @[Mux.scala 46:19:@11439.4]
  wire [7:0] _T_13626; // @[Mux.scala 46:16:@11440.4]
  wire  _T_13627; // @[Mux.scala 46:19:@11441.4]
  wire [7:0] _T_13628; // @[Mux.scala 46:16:@11442.4]
  wire  _T_13629; // @[Mux.scala 46:19:@11443.4]
  wire [7:0] _T_13630; // @[Mux.scala 46:16:@11444.4]
  wire  _T_13631; // @[Mux.scala 46:19:@11445.4]
  wire [7:0] _T_13632; // @[Mux.scala 46:16:@11446.4]
  wire  _T_13633; // @[Mux.scala 46:19:@11447.4]
  wire [7:0] _T_13634; // @[Mux.scala 46:16:@11448.4]
  wire  _T_13635; // @[Mux.scala 46:19:@11449.4]
  wire [7:0] _T_13636; // @[Mux.scala 46:16:@11450.4]
  wire  _T_13637; // @[Mux.scala 46:19:@11451.4]
  wire [7:0] _T_13638; // @[Mux.scala 46:16:@11452.4]
  wire  _T_13639; // @[Mux.scala 46:19:@11453.4]
  wire [7:0] _T_13640; // @[Mux.scala 46:16:@11454.4]
  wire  _T_13641; // @[Mux.scala 46:19:@11455.4]
  wire [7:0] _T_13642; // @[Mux.scala 46:16:@11456.4]
  wire  _T_13643; // @[Mux.scala 46:19:@11457.4]
  wire [7:0] _T_13644; // @[Mux.scala 46:16:@11458.4]
  wire  _T_13645; // @[Mux.scala 46:19:@11459.4]
  wire [7:0] _T_13646; // @[Mux.scala 46:16:@11460.4]
  wire  _T_13647; // @[Mux.scala 46:19:@11461.4]
  wire [7:0] _T_13648; // @[Mux.scala 46:16:@11462.4]
  wire  _T_13649; // @[Mux.scala 46:19:@11463.4]
  wire [7:0] _T_13650; // @[Mux.scala 46:16:@11464.4]
  wire  _T_13651; // @[Mux.scala 46:19:@11465.4]
  wire [7:0] _T_13652; // @[Mux.scala 46:16:@11466.4]
  wire  _T_13653; // @[Mux.scala 46:19:@11467.4]
  wire [7:0] _T_13654; // @[Mux.scala 46:16:@11468.4]
  wire  _T_13655; // @[Mux.scala 46:19:@11469.4]
  wire [7:0] _T_13656; // @[Mux.scala 46:16:@11470.4]
  wire  _T_13657; // @[Mux.scala 46:19:@11471.4]
  wire [7:0] _T_13658; // @[Mux.scala 46:16:@11472.4]
  wire  _T_13659; // @[Mux.scala 46:19:@11473.4]
  wire [7:0] _T_13660; // @[Mux.scala 46:16:@11474.4]
  wire  _T_13661; // @[Mux.scala 46:19:@11475.4]
  wire [7:0] _T_13662; // @[Mux.scala 46:16:@11476.4]
  wire  _T_13663; // @[Mux.scala 46:19:@11477.4]
  wire [7:0] _T_13664; // @[Mux.scala 46:16:@11478.4]
  wire  _T_13665; // @[Mux.scala 46:19:@11479.4]
  wire [7:0] _T_13666; // @[Mux.scala 46:16:@11480.4]
  wire  _T_13667; // @[Mux.scala 46:19:@11481.4]
  wire [7:0] _T_13668; // @[Mux.scala 46:16:@11482.4]
  wire  _T_13669; // @[Mux.scala 46:19:@11483.4]
  wire [7:0] _T_13670; // @[Mux.scala 46:16:@11484.4]
  wire  _T_13671; // @[Mux.scala 46:19:@11485.4]
  wire [7:0] _T_13672; // @[Mux.scala 46:16:@11486.4]
  wire  _T_13673; // @[Mux.scala 46:19:@11487.4]
  wire [7:0] _T_13674; // @[Mux.scala 46:16:@11488.4]
  wire  _T_13675; // @[Mux.scala 46:19:@11489.4]
  wire [7:0] _T_13676; // @[Mux.scala 46:16:@11490.4]
  wire  _T_13677; // @[Mux.scala 46:19:@11491.4]
  wire [7:0] _T_13678; // @[Mux.scala 46:16:@11492.4]
  wire  _T_13679; // @[Mux.scala 46:19:@11493.4]
  wire [7:0] _T_13680; // @[Mux.scala 46:16:@11494.4]
  wire  _T_13681; // @[Mux.scala 46:19:@11495.4]
  wire [7:0] _T_13682; // @[Mux.scala 46:16:@11496.4]
  wire  _T_13683; // @[Mux.scala 46:19:@11497.4]
  wire [7:0] _T_13684; // @[Mux.scala 46:16:@11498.4]
  wire  _T_13685; // @[Mux.scala 46:19:@11499.4]
  wire [7:0] _T_13686; // @[Mux.scala 46:16:@11500.4]
  wire  _T_13687; // @[Mux.scala 46:19:@11501.4]
  wire [7:0] _T_13688; // @[Mux.scala 46:16:@11502.4]
  wire  _T_13689; // @[Mux.scala 46:19:@11503.4]
  wire [7:0] _T_13690; // @[Mux.scala 46:16:@11504.4]
  wire  _T_13691; // @[Mux.scala 46:19:@11505.4]
  wire [7:0] _T_13692; // @[Mux.scala 46:16:@11506.4]
  wire  _T_13693; // @[Mux.scala 46:19:@11507.4]
  wire [7:0] _T_13694; // @[Mux.scala 46:16:@11508.4]
  wire  _T_13695; // @[Mux.scala 46:19:@11509.4]
  wire [7:0] _T_13696; // @[Mux.scala 46:16:@11510.4]
  wire  _T_13697; // @[Mux.scala 46:19:@11511.4]
  wire [7:0] _T_13698; // @[Mux.scala 46:16:@11512.4]
  wire  _T_13747; // @[Mux.scala 46:19:@11514.4]
  wire [7:0] _T_13748; // @[Mux.scala 46:16:@11515.4]
  wire  _T_13749; // @[Mux.scala 46:19:@11516.4]
  wire [7:0] _T_13750; // @[Mux.scala 46:16:@11517.4]
  wire  _T_13751; // @[Mux.scala 46:19:@11518.4]
  wire [7:0] _T_13752; // @[Mux.scala 46:16:@11519.4]
  wire  _T_13753; // @[Mux.scala 46:19:@11520.4]
  wire [7:0] _T_13754; // @[Mux.scala 46:16:@11521.4]
  wire  _T_13755; // @[Mux.scala 46:19:@11522.4]
  wire [7:0] _T_13756; // @[Mux.scala 46:16:@11523.4]
  wire  _T_13757; // @[Mux.scala 46:19:@11524.4]
  wire [7:0] _T_13758; // @[Mux.scala 46:16:@11525.4]
  wire  _T_13759; // @[Mux.scala 46:19:@11526.4]
  wire [7:0] _T_13760; // @[Mux.scala 46:16:@11527.4]
  wire  _T_13761; // @[Mux.scala 46:19:@11528.4]
  wire [7:0] _T_13762; // @[Mux.scala 46:16:@11529.4]
  wire  _T_13763; // @[Mux.scala 46:19:@11530.4]
  wire [7:0] _T_13764; // @[Mux.scala 46:16:@11531.4]
  wire  _T_13765; // @[Mux.scala 46:19:@11532.4]
  wire [7:0] _T_13766; // @[Mux.scala 46:16:@11533.4]
  wire  _T_13767; // @[Mux.scala 46:19:@11534.4]
  wire [7:0] _T_13768; // @[Mux.scala 46:16:@11535.4]
  wire  _T_13769; // @[Mux.scala 46:19:@11536.4]
  wire [7:0] _T_13770; // @[Mux.scala 46:16:@11537.4]
  wire  _T_13771; // @[Mux.scala 46:19:@11538.4]
  wire [7:0] _T_13772; // @[Mux.scala 46:16:@11539.4]
  wire  _T_13773; // @[Mux.scala 46:19:@11540.4]
  wire [7:0] _T_13774; // @[Mux.scala 46:16:@11541.4]
  wire  _T_13775; // @[Mux.scala 46:19:@11542.4]
  wire [7:0] _T_13776; // @[Mux.scala 46:16:@11543.4]
  wire  _T_13777; // @[Mux.scala 46:19:@11544.4]
  wire [7:0] _T_13778; // @[Mux.scala 46:16:@11545.4]
  wire  _T_13779; // @[Mux.scala 46:19:@11546.4]
  wire [7:0] _T_13780; // @[Mux.scala 46:16:@11547.4]
  wire  _T_13781; // @[Mux.scala 46:19:@11548.4]
  wire [7:0] _T_13782; // @[Mux.scala 46:16:@11549.4]
  wire  _T_13783; // @[Mux.scala 46:19:@11550.4]
  wire [7:0] _T_13784; // @[Mux.scala 46:16:@11551.4]
  wire  _T_13785; // @[Mux.scala 46:19:@11552.4]
  wire [7:0] _T_13786; // @[Mux.scala 46:16:@11553.4]
  wire  _T_13787; // @[Mux.scala 46:19:@11554.4]
  wire [7:0] _T_13788; // @[Mux.scala 46:16:@11555.4]
  wire  _T_13789; // @[Mux.scala 46:19:@11556.4]
  wire [7:0] _T_13790; // @[Mux.scala 46:16:@11557.4]
  wire  _T_13791; // @[Mux.scala 46:19:@11558.4]
  wire [7:0] _T_13792; // @[Mux.scala 46:16:@11559.4]
  wire  _T_13793; // @[Mux.scala 46:19:@11560.4]
  wire [7:0] _T_13794; // @[Mux.scala 46:16:@11561.4]
  wire  _T_13795; // @[Mux.scala 46:19:@11562.4]
  wire [7:0] _T_13796; // @[Mux.scala 46:16:@11563.4]
  wire  _T_13797; // @[Mux.scala 46:19:@11564.4]
  wire [7:0] _T_13798; // @[Mux.scala 46:16:@11565.4]
  wire  _T_13799; // @[Mux.scala 46:19:@11566.4]
  wire [7:0] _T_13800; // @[Mux.scala 46:16:@11567.4]
  wire  _T_13801; // @[Mux.scala 46:19:@11568.4]
  wire [7:0] _T_13802; // @[Mux.scala 46:16:@11569.4]
  wire  _T_13803; // @[Mux.scala 46:19:@11570.4]
  wire [7:0] _T_13804; // @[Mux.scala 46:16:@11571.4]
  wire  _T_13805; // @[Mux.scala 46:19:@11572.4]
  wire [7:0] _T_13806; // @[Mux.scala 46:16:@11573.4]
  wire  _T_13807; // @[Mux.scala 46:19:@11574.4]
  wire [7:0] _T_13808; // @[Mux.scala 46:16:@11575.4]
  wire  _T_13809; // @[Mux.scala 46:19:@11576.4]
  wire [7:0] _T_13810; // @[Mux.scala 46:16:@11577.4]
  wire  _T_13811; // @[Mux.scala 46:19:@11578.4]
  wire [7:0] _T_13812; // @[Mux.scala 46:16:@11579.4]
  wire  _T_13813; // @[Mux.scala 46:19:@11580.4]
  wire [7:0] _T_13814; // @[Mux.scala 46:16:@11581.4]
  wire  _T_13815; // @[Mux.scala 46:19:@11582.4]
  wire [7:0] _T_13816; // @[Mux.scala 46:16:@11583.4]
  wire  _T_13817; // @[Mux.scala 46:19:@11584.4]
  wire [7:0] _T_13818; // @[Mux.scala 46:16:@11585.4]
  wire  _T_13819; // @[Mux.scala 46:19:@11586.4]
  wire [7:0] _T_13820; // @[Mux.scala 46:16:@11587.4]
  wire  _T_13821; // @[Mux.scala 46:19:@11588.4]
  wire [7:0] _T_13822; // @[Mux.scala 46:16:@11589.4]
  wire  _T_13823; // @[Mux.scala 46:19:@11590.4]
  wire [7:0] _T_13824; // @[Mux.scala 46:16:@11591.4]
  wire  _T_13825; // @[Mux.scala 46:19:@11592.4]
  wire [7:0] _T_13826; // @[Mux.scala 46:16:@11593.4]
  wire  _T_13827; // @[Mux.scala 46:19:@11594.4]
  wire [7:0] _T_13828; // @[Mux.scala 46:16:@11595.4]
  wire  _T_13829; // @[Mux.scala 46:19:@11596.4]
  wire [7:0] _T_13830; // @[Mux.scala 46:16:@11597.4]
  wire  _T_13831; // @[Mux.scala 46:19:@11598.4]
  wire [7:0] _T_13832; // @[Mux.scala 46:16:@11599.4]
  wire  _T_13833; // @[Mux.scala 46:19:@11600.4]
  wire [7:0] _T_13834; // @[Mux.scala 46:16:@11601.4]
  wire  _T_13835; // @[Mux.scala 46:19:@11602.4]
  wire [7:0] _T_13836; // @[Mux.scala 46:16:@11603.4]
  wire  _T_13837; // @[Mux.scala 46:19:@11604.4]
  wire [7:0] _T_13838; // @[Mux.scala 46:16:@11605.4]
  wire  _T_13839; // @[Mux.scala 46:19:@11606.4]
  wire [7:0] _T_13840; // @[Mux.scala 46:16:@11607.4]
  wire  _T_13890; // @[Mux.scala 46:19:@11609.4]
  wire [7:0] _T_13891; // @[Mux.scala 46:16:@11610.4]
  wire  _T_13892; // @[Mux.scala 46:19:@11611.4]
  wire [7:0] _T_13893; // @[Mux.scala 46:16:@11612.4]
  wire  _T_13894; // @[Mux.scala 46:19:@11613.4]
  wire [7:0] _T_13895; // @[Mux.scala 46:16:@11614.4]
  wire  _T_13896; // @[Mux.scala 46:19:@11615.4]
  wire [7:0] _T_13897; // @[Mux.scala 46:16:@11616.4]
  wire  _T_13898; // @[Mux.scala 46:19:@11617.4]
  wire [7:0] _T_13899; // @[Mux.scala 46:16:@11618.4]
  wire  _T_13900; // @[Mux.scala 46:19:@11619.4]
  wire [7:0] _T_13901; // @[Mux.scala 46:16:@11620.4]
  wire  _T_13902; // @[Mux.scala 46:19:@11621.4]
  wire [7:0] _T_13903; // @[Mux.scala 46:16:@11622.4]
  wire  _T_13904; // @[Mux.scala 46:19:@11623.4]
  wire [7:0] _T_13905; // @[Mux.scala 46:16:@11624.4]
  wire  _T_13906; // @[Mux.scala 46:19:@11625.4]
  wire [7:0] _T_13907; // @[Mux.scala 46:16:@11626.4]
  wire  _T_13908; // @[Mux.scala 46:19:@11627.4]
  wire [7:0] _T_13909; // @[Mux.scala 46:16:@11628.4]
  wire  _T_13910; // @[Mux.scala 46:19:@11629.4]
  wire [7:0] _T_13911; // @[Mux.scala 46:16:@11630.4]
  wire  _T_13912; // @[Mux.scala 46:19:@11631.4]
  wire [7:0] _T_13913; // @[Mux.scala 46:16:@11632.4]
  wire  _T_13914; // @[Mux.scala 46:19:@11633.4]
  wire [7:0] _T_13915; // @[Mux.scala 46:16:@11634.4]
  wire  _T_13916; // @[Mux.scala 46:19:@11635.4]
  wire [7:0] _T_13917; // @[Mux.scala 46:16:@11636.4]
  wire  _T_13918; // @[Mux.scala 46:19:@11637.4]
  wire [7:0] _T_13919; // @[Mux.scala 46:16:@11638.4]
  wire  _T_13920; // @[Mux.scala 46:19:@11639.4]
  wire [7:0] _T_13921; // @[Mux.scala 46:16:@11640.4]
  wire  _T_13922; // @[Mux.scala 46:19:@11641.4]
  wire [7:0] _T_13923; // @[Mux.scala 46:16:@11642.4]
  wire  _T_13924; // @[Mux.scala 46:19:@11643.4]
  wire [7:0] _T_13925; // @[Mux.scala 46:16:@11644.4]
  wire  _T_13926; // @[Mux.scala 46:19:@11645.4]
  wire [7:0] _T_13927; // @[Mux.scala 46:16:@11646.4]
  wire  _T_13928; // @[Mux.scala 46:19:@11647.4]
  wire [7:0] _T_13929; // @[Mux.scala 46:16:@11648.4]
  wire  _T_13930; // @[Mux.scala 46:19:@11649.4]
  wire [7:0] _T_13931; // @[Mux.scala 46:16:@11650.4]
  wire  _T_13932; // @[Mux.scala 46:19:@11651.4]
  wire [7:0] _T_13933; // @[Mux.scala 46:16:@11652.4]
  wire  _T_13934; // @[Mux.scala 46:19:@11653.4]
  wire [7:0] _T_13935; // @[Mux.scala 46:16:@11654.4]
  wire  _T_13936; // @[Mux.scala 46:19:@11655.4]
  wire [7:0] _T_13937; // @[Mux.scala 46:16:@11656.4]
  wire  _T_13938; // @[Mux.scala 46:19:@11657.4]
  wire [7:0] _T_13939; // @[Mux.scala 46:16:@11658.4]
  wire  _T_13940; // @[Mux.scala 46:19:@11659.4]
  wire [7:0] _T_13941; // @[Mux.scala 46:16:@11660.4]
  wire  _T_13942; // @[Mux.scala 46:19:@11661.4]
  wire [7:0] _T_13943; // @[Mux.scala 46:16:@11662.4]
  wire  _T_13944; // @[Mux.scala 46:19:@11663.4]
  wire [7:0] _T_13945; // @[Mux.scala 46:16:@11664.4]
  wire  _T_13946; // @[Mux.scala 46:19:@11665.4]
  wire [7:0] _T_13947; // @[Mux.scala 46:16:@11666.4]
  wire  _T_13948; // @[Mux.scala 46:19:@11667.4]
  wire [7:0] _T_13949; // @[Mux.scala 46:16:@11668.4]
  wire  _T_13950; // @[Mux.scala 46:19:@11669.4]
  wire [7:0] _T_13951; // @[Mux.scala 46:16:@11670.4]
  wire  _T_13952; // @[Mux.scala 46:19:@11671.4]
  wire [7:0] _T_13953; // @[Mux.scala 46:16:@11672.4]
  wire  _T_13954; // @[Mux.scala 46:19:@11673.4]
  wire [7:0] _T_13955; // @[Mux.scala 46:16:@11674.4]
  wire  _T_13956; // @[Mux.scala 46:19:@11675.4]
  wire [7:0] _T_13957; // @[Mux.scala 46:16:@11676.4]
  wire  _T_13958; // @[Mux.scala 46:19:@11677.4]
  wire [7:0] _T_13959; // @[Mux.scala 46:16:@11678.4]
  wire  _T_13960; // @[Mux.scala 46:19:@11679.4]
  wire [7:0] _T_13961; // @[Mux.scala 46:16:@11680.4]
  wire  _T_13962; // @[Mux.scala 46:19:@11681.4]
  wire [7:0] _T_13963; // @[Mux.scala 46:16:@11682.4]
  wire  _T_13964; // @[Mux.scala 46:19:@11683.4]
  wire [7:0] _T_13965; // @[Mux.scala 46:16:@11684.4]
  wire  _T_13966; // @[Mux.scala 46:19:@11685.4]
  wire [7:0] _T_13967; // @[Mux.scala 46:16:@11686.4]
  wire  _T_13968; // @[Mux.scala 46:19:@11687.4]
  wire [7:0] _T_13969; // @[Mux.scala 46:16:@11688.4]
  wire  _T_13970; // @[Mux.scala 46:19:@11689.4]
  wire [7:0] _T_13971; // @[Mux.scala 46:16:@11690.4]
  wire  _T_13972; // @[Mux.scala 46:19:@11691.4]
  wire [7:0] _T_13973; // @[Mux.scala 46:16:@11692.4]
  wire  _T_13974; // @[Mux.scala 46:19:@11693.4]
  wire [7:0] _T_13975; // @[Mux.scala 46:16:@11694.4]
  wire  _T_13976; // @[Mux.scala 46:19:@11695.4]
  wire [7:0] _T_13977; // @[Mux.scala 46:16:@11696.4]
  wire  _T_13978; // @[Mux.scala 46:19:@11697.4]
  wire [7:0] _T_13979; // @[Mux.scala 46:16:@11698.4]
  wire  _T_13980; // @[Mux.scala 46:19:@11699.4]
  wire [7:0] _T_13981; // @[Mux.scala 46:16:@11700.4]
  wire  _T_13982; // @[Mux.scala 46:19:@11701.4]
  wire [7:0] _T_13983; // @[Mux.scala 46:16:@11702.4]
  wire  _T_13984; // @[Mux.scala 46:19:@11703.4]
  wire [7:0] _T_13985; // @[Mux.scala 46:16:@11704.4]
  wire  _T_14036; // @[Mux.scala 46:19:@11706.4]
  wire [7:0] _T_14037; // @[Mux.scala 46:16:@11707.4]
  wire  _T_14038; // @[Mux.scala 46:19:@11708.4]
  wire [7:0] _T_14039; // @[Mux.scala 46:16:@11709.4]
  wire  _T_14040; // @[Mux.scala 46:19:@11710.4]
  wire [7:0] _T_14041; // @[Mux.scala 46:16:@11711.4]
  wire  _T_14042; // @[Mux.scala 46:19:@11712.4]
  wire [7:0] _T_14043; // @[Mux.scala 46:16:@11713.4]
  wire  _T_14044; // @[Mux.scala 46:19:@11714.4]
  wire [7:0] _T_14045; // @[Mux.scala 46:16:@11715.4]
  wire  _T_14046; // @[Mux.scala 46:19:@11716.4]
  wire [7:0] _T_14047; // @[Mux.scala 46:16:@11717.4]
  wire  _T_14048; // @[Mux.scala 46:19:@11718.4]
  wire [7:0] _T_14049; // @[Mux.scala 46:16:@11719.4]
  wire  _T_14050; // @[Mux.scala 46:19:@11720.4]
  wire [7:0] _T_14051; // @[Mux.scala 46:16:@11721.4]
  wire  _T_14052; // @[Mux.scala 46:19:@11722.4]
  wire [7:0] _T_14053; // @[Mux.scala 46:16:@11723.4]
  wire  _T_14054; // @[Mux.scala 46:19:@11724.4]
  wire [7:0] _T_14055; // @[Mux.scala 46:16:@11725.4]
  wire  _T_14056; // @[Mux.scala 46:19:@11726.4]
  wire [7:0] _T_14057; // @[Mux.scala 46:16:@11727.4]
  wire  _T_14058; // @[Mux.scala 46:19:@11728.4]
  wire [7:0] _T_14059; // @[Mux.scala 46:16:@11729.4]
  wire  _T_14060; // @[Mux.scala 46:19:@11730.4]
  wire [7:0] _T_14061; // @[Mux.scala 46:16:@11731.4]
  wire  _T_14062; // @[Mux.scala 46:19:@11732.4]
  wire [7:0] _T_14063; // @[Mux.scala 46:16:@11733.4]
  wire  _T_14064; // @[Mux.scala 46:19:@11734.4]
  wire [7:0] _T_14065; // @[Mux.scala 46:16:@11735.4]
  wire  _T_14066; // @[Mux.scala 46:19:@11736.4]
  wire [7:0] _T_14067; // @[Mux.scala 46:16:@11737.4]
  wire  _T_14068; // @[Mux.scala 46:19:@11738.4]
  wire [7:0] _T_14069; // @[Mux.scala 46:16:@11739.4]
  wire  _T_14070; // @[Mux.scala 46:19:@11740.4]
  wire [7:0] _T_14071; // @[Mux.scala 46:16:@11741.4]
  wire  _T_14072; // @[Mux.scala 46:19:@11742.4]
  wire [7:0] _T_14073; // @[Mux.scala 46:16:@11743.4]
  wire  _T_14074; // @[Mux.scala 46:19:@11744.4]
  wire [7:0] _T_14075; // @[Mux.scala 46:16:@11745.4]
  wire  _T_14076; // @[Mux.scala 46:19:@11746.4]
  wire [7:0] _T_14077; // @[Mux.scala 46:16:@11747.4]
  wire  _T_14078; // @[Mux.scala 46:19:@11748.4]
  wire [7:0] _T_14079; // @[Mux.scala 46:16:@11749.4]
  wire  _T_14080; // @[Mux.scala 46:19:@11750.4]
  wire [7:0] _T_14081; // @[Mux.scala 46:16:@11751.4]
  wire  _T_14082; // @[Mux.scala 46:19:@11752.4]
  wire [7:0] _T_14083; // @[Mux.scala 46:16:@11753.4]
  wire  _T_14084; // @[Mux.scala 46:19:@11754.4]
  wire [7:0] _T_14085; // @[Mux.scala 46:16:@11755.4]
  wire  _T_14086; // @[Mux.scala 46:19:@11756.4]
  wire [7:0] _T_14087; // @[Mux.scala 46:16:@11757.4]
  wire  _T_14088; // @[Mux.scala 46:19:@11758.4]
  wire [7:0] _T_14089; // @[Mux.scala 46:16:@11759.4]
  wire  _T_14090; // @[Mux.scala 46:19:@11760.4]
  wire [7:0] _T_14091; // @[Mux.scala 46:16:@11761.4]
  wire  _T_14092; // @[Mux.scala 46:19:@11762.4]
  wire [7:0] _T_14093; // @[Mux.scala 46:16:@11763.4]
  wire  _T_14094; // @[Mux.scala 46:19:@11764.4]
  wire [7:0] _T_14095; // @[Mux.scala 46:16:@11765.4]
  wire  _T_14096; // @[Mux.scala 46:19:@11766.4]
  wire [7:0] _T_14097; // @[Mux.scala 46:16:@11767.4]
  wire  _T_14098; // @[Mux.scala 46:19:@11768.4]
  wire [7:0] _T_14099; // @[Mux.scala 46:16:@11769.4]
  wire  _T_14100; // @[Mux.scala 46:19:@11770.4]
  wire [7:0] _T_14101; // @[Mux.scala 46:16:@11771.4]
  wire  _T_14102; // @[Mux.scala 46:19:@11772.4]
  wire [7:0] _T_14103; // @[Mux.scala 46:16:@11773.4]
  wire  _T_14104; // @[Mux.scala 46:19:@11774.4]
  wire [7:0] _T_14105; // @[Mux.scala 46:16:@11775.4]
  wire  _T_14106; // @[Mux.scala 46:19:@11776.4]
  wire [7:0] _T_14107; // @[Mux.scala 46:16:@11777.4]
  wire  _T_14108; // @[Mux.scala 46:19:@11778.4]
  wire [7:0] _T_14109; // @[Mux.scala 46:16:@11779.4]
  wire  _T_14110; // @[Mux.scala 46:19:@11780.4]
  wire [7:0] _T_14111; // @[Mux.scala 46:16:@11781.4]
  wire  _T_14112; // @[Mux.scala 46:19:@11782.4]
  wire [7:0] _T_14113; // @[Mux.scala 46:16:@11783.4]
  wire  _T_14114; // @[Mux.scala 46:19:@11784.4]
  wire [7:0] _T_14115; // @[Mux.scala 46:16:@11785.4]
  wire  _T_14116; // @[Mux.scala 46:19:@11786.4]
  wire [7:0] _T_14117; // @[Mux.scala 46:16:@11787.4]
  wire  _T_14118; // @[Mux.scala 46:19:@11788.4]
  wire [7:0] _T_14119; // @[Mux.scala 46:16:@11789.4]
  wire  _T_14120; // @[Mux.scala 46:19:@11790.4]
  wire [7:0] _T_14121; // @[Mux.scala 46:16:@11791.4]
  wire  _T_14122; // @[Mux.scala 46:19:@11792.4]
  wire [7:0] _T_14123; // @[Mux.scala 46:16:@11793.4]
  wire  _T_14124; // @[Mux.scala 46:19:@11794.4]
  wire [7:0] _T_14125; // @[Mux.scala 46:16:@11795.4]
  wire  _T_14126; // @[Mux.scala 46:19:@11796.4]
  wire [7:0] _T_14127; // @[Mux.scala 46:16:@11797.4]
  wire  _T_14128; // @[Mux.scala 46:19:@11798.4]
  wire [7:0] _T_14129; // @[Mux.scala 46:16:@11799.4]
  wire  _T_14130; // @[Mux.scala 46:19:@11800.4]
  wire [7:0] _T_14131; // @[Mux.scala 46:16:@11801.4]
  wire  _T_14132; // @[Mux.scala 46:19:@11802.4]
  wire [7:0] _T_14133; // @[Mux.scala 46:16:@11803.4]
  wire  _T_14185; // @[Mux.scala 46:19:@11805.4]
  wire [7:0] _T_14186; // @[Mux.scala 46:16:@11806.4]
  wire  _T_14187; // @[Mux.scala 46:19:@11807.4]
  wire [7:0] _T_14188; // @[Mux.scala 46:16:@11808.4]
  wire  _T_14189; // @[Mux.scala 46:19:@11809.4]
  wire [7:0] _T_14190; // @[Mux.scala 46:16:@11810.4]
  wire  _T_14191; // @[Mux.scala 46:19:@11811.4]
  wire [7:0] _T_14192; // @[Mux.scala 46:16:@11812.4]
  wire  _T_14193; // @[Mux.scala 46:19:@11813.4]
  wire [7:0] _T_14194; // @[Mux.scala 46:16:@11814.4]
  wire  _T_14195; // @[Mux.scala 46:19:@11815.4]
  wire [7:0] _T_14196; // @[Mux.scala 46:16:@11816.4]
  wire  _T_14197; // @[Mux.scala 46:19:@11817.4]
  wire [7:0] _T_14198; // @[Mux.scala 46:16:@11818.4]
  wire  _T_14199; // @[Mux.scala 46:19:@11819.4]
  wire [7:0] _T_14200; // @[Mux.scala 46:16:@11820.4]
  wire  _T_14201; // @[Mux.scala 46:19:@11821.4]
  wire [7:0] _T_14202; // @[Mux.scala 46:16:@11822.4]
  wire  _T_14203; // @[Mux.scala 46:19:@11823.4]
  wire [7:0] _T_14204; // @[Mux.scala 46:16:@11824.4]
  wire  _T_14205; // @[Mux.scala 46:19:@11825.4]
  wire [7:0] _T_14206; // @[Mux.scala 46:16:@11826.4]
  wire  _T_14207; // @[Mux.scala 46:19:@11827.4]
  wire [7:0] _T_14208; // @[Mux.scala 46:16:@11828.4]
  wire  _T_14209; // @[Mux.scala 46:19:@11829.4]
  wire [7:0] _T_14210; // @[Mux.scala 46:16:@11830.4]
  wire  _T_14211; // @[Mux.scala 46:19:@11831.4]
  wire [7:0] _T_14212; // @[Mux.scala 46:16:@11832.4]
  wire  _T_14213; // @[Mux.scala 46:19:@11833.4]
  wire [7:0] _T_14214; // @[Mux.scala 46:16:@11834.4]
  wire  _T_14215; // @[Mux.scala 46:19:@11835.4]
  wire [7:0] _T_14216; // @[Mux.scala 46:16:@11836.4]
  wire  _T_14217; // @[Mux.scala 46:19:@11837.4]
  wire [7:0] _T_14218; // @[Mux.scala 46:16:@11838.4]
  wire  _T_14219; // @[Mux.scala 46:19:@11839.4]
  wire [7:0] _T_14220; // @[Mux.scala 46:16:@11840.4]
  wire  _T_14221; // @[Mux.scala 46:19:@11841.4]
  wire [7:0] _T_14222; // @[Mux.scala 46:16:@11842.4]
  wire  _T_14223; // @[Mux.scala 46:19:@11843.4]
  wire [7:0] _T_14224; // @[Mux.scala 46:16:@11844.4]
  wire  _T_14225; // @[Mux.scala 46:19:@11845.4]
  wire [7:0] _T_14226; // @[Mux.scala 46:16:@11846.4]
  wire  _T_14227; // @[Mux.scala 46:19:@11847.4]
  wire [7:0] _T_14228; // @[Mux.scala 46:16:@11848.4]
  wire  _T_14229; // @[Mux.scala 46:19:@11849.4]
  wire [7:0] _T_14230; // @[Mux.scala 46:16:@11850.4]
  wire  _T_14231; // @[Mux.scala 46:19:@11851.4]
  wire [7:0] _T_14232; // @[Mux.scala 46:16:@11852.4]
  wire  _T_14233; // @[Mux.scala 46:19:@11853.4]
  wire [7:0] _T_14234; // @[Mux.scala 46:16:@11854.4]
  wire  _T_14235; // @[Mux.scala 46:19:@11855.4]
  wire [7:0] _T_14236; // @[Mux.scala 46:16:@11856.4]
  wire  _T_14237; // @[Mux.scala 46:19:@11857.4]
  wire [7:0] _T_14238; // @[Mux.scala 46:16:@11858.4]
  wire  _T_14239; // @[Mux.scala 46:19:@11859.4]
  wire [7:0] _T_14240; // @[Mux.scala 46:16:@11860.4]
  wire  _T_14241; // @[Mux.scala 46:19:@11861.4]
  wire [7:0] _T_14242; // @[Mux.scala 46:16:@11862.4]
  wire  _T_14243; // @[Mux.scala 46:19:@11863.4]
  wire [7:0] _T_14244; // @[Mux.scala 46:16:@11864.4]
  wire  _T_14245; // @[Mux.scala 46:19:@11865.4]
  wire [7:0] _T_14246; // @[Mux.scala 46:16:@11866.4]
  wire  _T_14247; // @[Mux.scala 46:19:@11867.4]
  wire [7:0] _T_14248; // @[Mux.scala 46:16:@11868.4]
  wire  _T_14249; // @[Mux.scala 46:19:@11869.4]
  wire [7:0] _T_14250; // @[Mux.scala 46:16:@11870.4]
  wire  _T_14251; // @[Mux.scala 46:19:@11871.4]
  wire [7:0] _T_14252; // @[Mux.scala 46:16:@11872.4]
  wire  _T_14253; // @[Mux.scala 46:19:@11873.4]
  wire [7:0] _T_14254; // @[Mux.scala 46:16:@11874.4]
  wire  _T_14255; // @[Mux.scala 46:19:@11875.4]
  wire [7:0] _T_14256; // @[Mux.scala 46:16:@11876.4]
  wire  _T_14257; // @[Mux.scala 46:19:@11877.4]
  wire [7:0] _T_14258; // @[Mux.scala 46:16:@11878.4]
  wire  _T_14259; // @[Mux.scala 46:19:@11879.4]
  wire [7:0] _T_14260; // @[Mux.scala 46:16:@11880.4]
  wire  _T_14261; // @[Mux.scala 46:19:@11881.4]
  wire [7:0] _T_14262; // @[Mux.scala 46:16:@11882.4]
  wire  _T_14263; // @[Mux.scala 46:19:@11883.4]
  wire [7:0] _T_14264; // @[Mux.scala 46:16:@11884.4]
  wire  _T_14265; // @[Mux.scala 46:19:@11885.4]
  wire [7:0] _T_14266; // @[Mux.scala 46:16:@11886.4]
  wire  _T_14267; // @[Mux.scala 46:19:@11887.4]
  wire [7:0] _T_14268; // @[Mux.scala 46:16:@11888.4]
  wire  _T_14269; // @[Mux.scala 46:19:@11889.4]
  wire [7:0] _T_14270; // @[Mux.scala 46:16:@11890.4]
  wire  _T_14271; // @[Mux.scala 46:19:@11891.4]
  wire [7:0] _T_14272; // @[Mux.scala 46:16:@11892.4]
  wire  _T_14273; // @[Mux.scala 46:19:@11893.4]
  wire [7:0] _T_14274; // @[Mux.scala 46:16:@11894.4]
  wire  _T_14275; // @[Mux.scala 46:19:@11895.4]
  wire [7:0] _T_14276; // @[Mux.scala 46:16:@11896.4]
  wire  _T_14277; // @[Mux.scala 46:19:@11897.4]
  wire [7:0] _T_14278; // @[Mux.scala 46:16:@11898.4]
  wire  _T_14279; // @[Mux.scala 46:19:@11899.4]
  wire [7:0] _T_14280; // @[Mux.scala 46:16:@11900.4]
  wire  _T_14281; // @[Mux.scala 46:19:@11901.4]
  wire [7:0] _T_14282; // @[Mux.scala 46:16:@11902.4]
  wire  _T_14283; // @[Mux.scala 46:19:@11903.4]
  wire [7:0] _T_14284; // @[Mux.scala 46:16:@11904.4]
  wire  _T_14337; // @[Mux.scala 46:19:@11906.4]
  wire [7:0] _T_14338; // @[Mux.scala 46:16:@11907.4]
  wire  _T_14339; // @[Mux.scala 46:19:@11908.4]
  wire [7:0] _T_14340; // @[Mux.scala 46:16:@11909.4]
  wire  _T_14341; // @[Mux.scala 46:19:@11910.4]
  wire [7:0] _T_14342; // @[Mux.scala 46:16:@11911.4]
  wire  _T_14343; // @[Mux.scala 46:19:@11912.4]
  wire [7:0] _T_14344; // @[Mux.scala 46:16:@11913.4]
  wire  _T_14345; // @[Mux.scala 46:19:@11914.4]
  wire [7:0] _T_14346; // @[Mux.scala 46:16:@11915.4]
  wire  _T_14347; // @[Mux.scala 46:19:@11916.4]
  wire [7:0] _T_14348; // @[Mux.scala 46:16:@11917.4]
  wire  _T_14349; // @[Mux.scala 46:19:@11918.4]
  wire [7:0] _T_14350; // @[Mux.scala 46:16:@11919.4]
  wire  _T_14351; // @[Mux.scala 46:19:@11920.4]
  wire [7:0] _T_14352; // @[Mux.scala 46:16:@11921.4]
  wire  _T_14353; // @[Mux.scala 46:19:@11922.4]
  wire [7:0] _T_14354; // @[Mux.scala 46:16:@11923.4]
  wire  _T_14355; // @[Mux.scala 46:19:@11924.4]
  wire [7:0] _T_14356; // @[Mux.scala 46:16:@11925.4]
  wire  _T_14357; // @[Mux.scala 46:19:@11926.4]
  wire [7:0] _T_14358; // @[Mux.scala 46:16:@11927.4]
  wire  _T_14359; // @[Mux.scala 46:19:@11928.4]
  wire [7:0] _T_14360; // @[Mux.scala 46:16:@11929.4]
  wire  _T_14361; // @[Mux.scala 46:19:@11930.4]
  wire [7:0] _T_14362; // @[Mux.scala 46:16:@11931.4]
  wire  _T_14363; // @[Mux.scala 46:19:@11932.4]
  wire [7:0] _T_14364; // @[Mux.scala 46:16:@11933.4]
  wire  _T_14365; // @[Mux.scala 46:19:@11934.4]
  wire [7:0] _T_14366; // @[Mux.scala 46:16:@11935.4]
  wire  _T_14367; // @[Mux.scala 46:19:@11936.4]
  wire [7:0] _T_14368; // @[Mux.scala 46:16:@11937.4]
  wire  _T_14369; // @[Mux.scala 46:19:@11938.4]
  wire [7:0] _T_14370; // @[Mux.scala 46:16:@11939.4]
  wire  _T_14371; // @[Mux.scala 46:19:@11940.4]
  wire [7:0] _T_14372; // @[Mux.scala 46:16:@11941.4]
  wire  _T_14373; // @[Mux.scala 46:19:@11942.4]
  wire [7:0] _T_14374; // @[Mux.scala 46:16:@11943.4]
  wire  _T_14375; // @[Mux.scala 46:19:@11944.4]
  wire [7:0] _T_14376; // @[Mux.scala 46:16:@11945.4]
  wire  _T_14377; // @[Mux.scala 46:19:@11946.4]
  wire [7:0] _T_14378; // @[Mux.scala 46:16:@11947.4]
  wire  _T_14379; // @[Mux.scala 46:19:@11948.4]
  wire [7:0] _T_14380; // @[Mux.scala 46:16:@11949.4]
  wire  _T_14381; // @[Mux.scala 46:19:@11950.4]
  wire [7:0] _T_14382; // @[Mux.scala 46:16:@11951.4]
  wire  _T_14383; // @[Mux.scala 46:19:@11952.4]
  wire [7:0] _T_14384; // @[Mux.scala 46:16:@11953.4]
  wire  _T_14385; // @[Mux.scala 46:19:@11954.4]
  wire [7:0] _T_14386; // @[Mux.scala 46:16:@11955.4]
  wire  _T_14387; // @[Mux.scala 46:19:@11956.4]
  wire [7:0] _T_14388; // @[Mux.scala 46:16:@11957.4]
  wire  _T_14389; // @[Mux.scala 46:19:@11958.4]
  wire [7:0] _T_14390; // @[Mux.scala 46:16:@11959.4]
  wire  _T_14391; // @[Mux.scala 46:19:@11960.4]
  wire [7:0] _T_14392; // @[Mux.scala 46:16:@11961.4]
  wire  _T_14393; // @[Mux.scala 46:19:@11962.4]
  wire [7:0] _T_14394; // @[Mux.scala 46:16:@11963.4]
  wire  _T_14395; // @[Mux.scala 46:19:@11964.4]
  wire [7:0] _T_14396; // @[Mux.scala 46:16:@11965.4]
  wire  _T_14397; // @[Mux.scala 46:19:@11966.4]
  wire [7:0] _T_14398; // @[Mux.scala 46:16:@11967.4]
  wire  _T_14399; // @[Mux.scala 46:19:@11968.4]
  wire [7:0] _T_14400; // @[Mux.scala 46:16:@11969.4]
  wire  _T_14401; // @[Mux.scala 46:19:@11970.4]
  wire [7:0] _T_14402; // @[Mux.scala 46:16:@11971.4]
  wire  _T_14403; // @[Mux.scala 46:19:@11972.4]
  wire [7:0] _T_14404; // @[Mux.scala 46:16:@11973.4]
  wire  _T_14405; // @[Mux.scala 46:19:@11974.4]
  wire [7:0] _T_14406; // @[Mux.scala 46:16:@11975.4]
  wire  _T_14407; // @[Mux.scala 46:19:@11976.4]
  wire [7:0] _T_14408; // @[Mux.scala 46:16:@11977.4]
  wire  _T_14409; // @[Mux.scala 46:19:@11978.4]
  wire [7:0] _T_14410; // @[Mux.scala 46:16:@11979.4]
  wire  _T_14411; // @[Mux.scala 46:19:@11980.4]
  wire [7:0] _T_14412; // @[Mux.scala 46:16:@11981.4]
  wire  _T_14413; // @[Mux.scala 46:19:@11982.4]
  wire [7:0] _T_14414; // @[Mux.scala 46:16:@11983.4]
  wire  _T_14415; // @[Mux.scala 46:19:@11984.4]
  wire [7:0] _T_14416; // @[Mux.scala 46:16:@11985.4]
  wire  _T_14417; // @[Mux.scala 46:19:@11986.4]
  wire [7:0] _T_14418; // @[Mux.scala 46:16:@11987.4]
  wire  _T_14419; // @[Mux.scala 46:19:@11988.4]
  wire [7:0] _T_14420; // @[Mux.scala 46:16:@11989.4]
  wire  _T_14421; // @[Mux.scala 46:19:@11990.4]
  wire [7:0] _T_14422; // @[Mux.scala 46:16:@11991.4]
  wire  _T_14423; // @[Mux.scala 46:19:@11992.4]
  wire [7:0] _T_14424; // @[Mux.scala 46:16:@11993.4]
  wire  _T_14425; // @[Mux.scala 46:19:@11994.4]
  wire [7:0] _T_14426; // @[Mux.scala 46:16:@11995.4]
  wire  _T_14427; // @[Mux.scala 46:19:@11996.4]
  wire [7:0] _T_14428; // @[Mux.scala 46:16:@11997.4]
  wire  _T_14429; // @[Mux.scala 46:19:@11998.4]
  wire [7:0] _T_14430; // @[Mux.scala 46:16:@11999.4]
  wire  _T_14431; // @[Mux.scala 46:19:@12000.4]
  wire [7:0] _T_14432; // @[Mux.scala 46:16:@12001.4]
  wire  _T_14433; // @[Mux.scala 46:19:@12002.4]
  wire [7:0] _T_14434; // @[Mux.scala 46:16:@12003.4]
  wire  _T_14435; // @[Mux.scala 46:19:@12004.4]
  wire [7:0] _T_14436; // @[Mux.scala 46:16:@12005.4]
  wire  _T_14437; // @[Mux.scala 46:19:@12006.4]
  wire [7:0] _T_14438; // @[Mux.scala 46:16:@12007.4]
  wire  _T_14492; // @[Mux.scala 46:19:@12009.4]
  wire [7:0] _T_14493; // @[Mux.scala 46:16:@12010.4]
  wire  _T_14494; // @[Mux.scala 46:19:@12011.4]
  wire [7:0] _T_14495; // @[Mux.scala 46:16:@12012.4]
  wire  _T_14496; // @[Mux.scala 46:19:@12013.4]
  wire [7:0] _T_14497; // @[Mux.scala 46:16:@12014.4]
  wire  _T_14498; // @[Mux.scala 46:19:@12015.4]
  wire [7:0] _T_14499; // @[Mux.scala 46:16:@12016.4]
  wire  _T_14500; // @[Mux.scala 46:19:@12017.4]
  wire [7:0] _T_14501; // @[Mux.scala 46:16:@12018.4]
  wire  _T_14502; // @[Mux.scala 46:19:@12019.4]
  wire [7:0] _T_14503; // @[Mux.scala 46:16:@12020.4]
  wire  _T_14504; // @[Mux.scala 46:19:@12021.4]
  wire [7:0] _T_14505; // @[Mux.scala 46:16:@12022.4]
  wire  _T_14506; // @[Mux.scala 46:19:@12023.4]
  wire [7:0] _T_14507; // @[Mux.scala 46:16:@12024.4]
  wire  _T_14508; // @[Mux.scala 46:19:@12025.4]
  wire [7:0] _T_14509; // @[Mux.scala 46:16:@12026.4]
  wire  _T_14510; // @[Mux.scala 46:19:@12027.4]
  wire [7:0] _T_14511; // @[Mux.scala 46:16:@12028.4]
  wire  _T_14512; // @[Mux.scala 46:19:@12029.4]
  wire [7:0] _T_14513; // @[Mux.scala 46:16:@12030.4]
  wire  _T_14514; // @[Mux.scala 46:19:@12031.4]
  wire [7:0] _T_14515; // @[Mux.scala 46:16:@12032.4]
  wire  _T_14516; // @[Mux.scala 46:19:@12033.4]
  wire [7:0] _T_14517; // @[Mux.scala 46:16:@12034.4]
  wire  _T_14518; // @[Mux.scala 46:19:@12035.4]
  wire [7:0] _T_14519; // @[Mux.scala 46:16:@12036.4]
  wire  _T_14520; // @[Mux.scala 46:19:@12037.4]
  wire [7:0] _T_14521; // @[Mux.scala 46:16:@12038.4]
  wire  _T_14522; // @[Mux.scala 46:19:@12039.4]
  wire [7:0] _T_14523; // @[Mux.scala 46:16:@12040.4]
  wire  _T_14524; // @[Mux.scala 46:19:@12041.4]
  wire [7:0] _T_14525; // @[Mux.scala 46:16:@12042.4]
  wire  _T_14526; // @[Mux.scala 46:19:@12043.4]
  wire [7:0] _T_14527; // @[Mux.scala 46:16:@12044.4]
  wire  _T_14528; // @[Mux.scala 46:19:@12045.4]
  wire [7:0] _T_14529; // @[Mux.scala 46:16:@12046.4]
  wire  _T_14530; // @[Mux.scala 46:19:@12047.4]
  wire [7:0] _T_14531; // @[Mux.scala 46:16:@12048.4]
  wire  _T_14532; // @[Mux.scala 46:19:@12049.4]
  wire [7:0] _T_14533; // @[Mux.scala 46:16:@12050.4]
  wire  _T_14534; // @[Mux.scala 46:19:@12051.4]
  wire [7:0] _T_14535; // @[Mux.scala 46:16:@12052.4]
  wire  _T_14536; // @[Mux.scala 46:19:@12053.4]
  wire [7:0] _T_14537; // @[Mux.scala 46:16:@12054.4]
  wire  _T_14538; // @[Mux.scala 46:19:@12055.4]
  wire [7:0] _T_14539; // @[Mux.scala 46:16:@12056.4]
  wire  _T_14540; // @[Mux.scala 46:19:@12057.4]
  wire [7:0] _T_14541; // @[Mux.scala 46:16:@12058.4]
  wire  _T_14542; // @[Mux.scala 46:19:@12059.4]
  wire [7:0] _T_14543; // @[Mux.scala 46:16:@12060.4]
  wire  _T_14544; // @[Mux.scala 46:19:@12061.4]
  wire [7:0] _T_14545; // @[Mux.scala 46:16:@12062.4]
  wire  _T_14546; // @[Mux.scala 46:19:@12063.4]
  wire [7:0] _T_14547; // @[Mux.scala 46:16:@12064.4]
  wire  _T_14548; // @[Mux.scala 46:19:@12065.4]
  wire [7:0] _T_14549; // @[Mux.scala 46:16:@12066.4]
  wire  _T_14550; // @[Mux.scala 46:19:@12067.4]
  wire [7:0] _T_14551; // @[Mux.scala 46:16:@12068.4]
  wire  _T_14552; // @[Mux.scala 46:19:@12069.4]
  wire [7:0] _T_14553; // @[Mux.scala 46:16:@12070.4]
  wire  _T_14554; // @[Mux.scala 46:19:@12071.4]
  wire [7:0] _T_14555; // @[Mux.scala 46:16:@12072.4]
  wire  _T_14556; // @[Mux.scala 46:19:@12073.4]
  wire [7:0] _T_14557; // @[Mux.scala 46:16:@12074.4]
  wire  _T_14558; // @[Mux.scala 46:19:@12075.4]
  wire [7:0] _T_14559; // @[Mux.scala 46:16:@12076.4]
  wire  _T_14560; // @[Mux.scala 46:19:@12077.4]
  wire [7:0] _T_14561; // @[Mux.scala 46:16:@12078.4]
  wire  _T_14562; // @[Mux.scala 46:19:@12079.4]
  wire [7:0] _T_14563; // @[Mux.scala 46:16:@12080.4]
  wire  _T_14564; // @[Mux.scala 46:19:@12081.4]
  wire [7:0] _T_14565; // @[Mux.scala 46:16:@12082.4]
  wire  _T_14566; // @[Mux.scala 46:19:@12083.4]
  wire [7:0] _T_14567; // @[Mux.scala 46:16:@12084.4]
  wire  _T_14568; // @[Mux.scala 46:19:@12085.4]
  wire [7:0] _T_14569; // @[Mux.scala 46:16:@12086.4]
  wire  _T_14570; // @[Mux.scala 46:19:@12087.4]
  wire [7:0] _T_14571; // @[Mux.scala 46:16:@12088.4]
  wire  _T_14572; // @[Mux.scala 46:19:@12089.4]
  wire [7:0] _T_14573; // @[Mux.scala 46:16:@12090.4]
  wire  _T_14574; // @[Mux.scala 46:19:@12091.4]
  wire [7:0] _T_14575; // @[Mux.scala 46:16:@12092.4]
  wire  _T_14576; // @[Mux.scala 46:19:@12093.4]
  wire [7:0] _T_14577; // @[Mux.scala 46:16:@12094.4]
  wire  _T_14578; // @[Mux.scala 46:19:@12095.4]
  wire [7:0] _T_14579; // @[Mux.scala 46:16:@12096.4]
  wire  _T_14580; // @[Mux.scala 46:19:@12097.4]
  wire [7:0] _T_14581; // @[Mux.scala 46:16:@12098.4]
  wire  _T_14582; // @[Mux.scala 46:19:@12099.4]
  wire [7:0] _T_14583; // @[Mux.scala 46:16:@12100.4]
  wire  _T_14584; // @[Mux.scala 46:19:@12101.4]
  wire [7:0] _T_14585; // @[Mux.scala 46:16:@12102.4]
  wire  _T_14586; // @[Mux.scala 46:19:@12103.4]
  wire [7:0] _T_14587; // @[Mux.scala 46:16:@12104.4]
  wire  _T_14588; // @[Mux.scala 46:19:@12105.4]
  wire [7:0] _T_14589; // @[Mux.scala 46:16:@12106.4]
  wire  _T_14590; // @[Mux.scala 46:19:@12107.4]
  wire [7:0] _T_14591; // @[Mux.scala 46:16:@12108.4]
  wire  _T_14592; // @[Mux.scala 46:19:@12109.4]
  wire [7:0] _T_14593; // @[Mux.scala 46:16:@12110.4]
  wire  _T_14594; // @[Mux.scala 46:19:@12111.4]
  wire [7:0] _T_14595; // @[Mux.scala 46:16:@12112.4]
  wire  _T_14650; // @[Mux.scala 46:19:@12114.4]
  wire [7:0] _T_14651; // @[Mux.scala 46:16:@12115.4]
  wire  _T_14652; // @[Mux.scala 46:19:@12116.4]
  wire [7:0] _T_14653; // @[Mux.scala 46:16:@12117.4]
  wire  _T_14654; // @[Mux.scala 46:19:@12118.4]
  wire [7:0] _T_14655; // @[Mux.scala 46:16:@12119.4]
  wire  _T_14656; // @[Mux.scala 46:19:@12120.4]
  wire [7:0] _T_14657; // @[Mux.scala 46:16:@12121.4]
  wire  _T_14658; // @[Mux.scala 46:19:@12122.4]
  wire [7:0] _T_14659; // @[Mux.scala 46:16:@12123.4]
  wire  _T_14660; // @[Mux.scala 46:19:@12124.4]
  wire [7:0] _T_14661; // @[Mux.scala 46:16:@12125.4]
  wire  _T_14662; // @[Mux.scala 46:19:@12126.4]
  wire [7:0] _T_14663; // @[Mux.scala 46:16:@12127.4]
  wire  _T_14664; // @[Mux.scala 46:19:@12128.4]
  wire [7:0] _T_14665; // @[Mux.scala 46:16:@12129.4]
  wire  _T_14666; // @[Mux.scala 46:19:@12130.4]
  wire [7:0] _T_14667; // @[Mux.scala 46:16:@12131.4]
  wire  _T_14668; // @[Mux.scala 46:19:@12132.4]
  wire [7:0] _T_14669; // @[Mux.scala 46:16:@12133.4]
  wire  _T_14670; // @[Mux.scala 46:19:@12134.4]
  wire [7:0] _T_14671; // @[Mux.scala 46:16:@12135.4]
  wire  _T_14672; // @[Mux.scala 46:19:@12136.4]
  wire [7:0] _T_14673; // @[Mux.scala 46:16:@12137.4]
  wire  _T_14674; // @[Mux.scala 46:19:@12138.4]
  wire [7:0] _T_14675; // @[Mux.scala 46:16:@12139.4]
  wire  _T_14676; // @[Mux.scala 46:19:@12140.4]
  wire [7:0] _T_14677; // @[Mux.scala 46:16:@12141.4]
  wire  _T_14678; // @[Mux.scala 46:19:@12142.4]
  wire [7:0] _T_14679; // @[Mux.scala 46:16:@12143.4]
  wire  _T_14680; // @[Mux.scala 46:19:@12144.4]
  wire [7:0] _T_14681; // @[Mux.scala 46:16:@12145.4]
  wire  _T_14682; // @[Mux.scala 46:19:@12146.4]
  wire [7:0] _T_14683; // @[Mux.scala 46:16:@12147.4]
  wire  _T_14684; // @[Mux.scala 46:19:@12148.4]
  wire [7:0] _T_14685; // @[Mux.scala 46:16:@12149.4]
  wire  _T_14686; // @[Mux.scala 46:19:@12150.4]
  wire [7:0] _T_14687; // @[Mux.scala 46:16:@12151.4]
  wire  _T_14688; // @[Mux.scala 46:19:@12152.4]
  wire [7:0] _T_14689; // @[Mux.scala 46:16:@12153.4]
  wire  _T_14690; // @[Mux.scala 46:19:@12154.4]
  wire [7:0] _T_14691; // @[Mux.scala 46:16:@12155.4]
  wire  _T_14692; // @[Mux.scala 46:19:@12156.4]
  wire [7:0] _T_14693; // @[Mux.scala 46:16:@12157.4]
  wire  _T_14694; // @[Mux.scala 46:19:@12158.4]
  wire [7:0] _T_14695; // @[Mux.scala 46:16:@12159.4]
  wire  _T_14696; // @[Mux.scala 46:19:@12160.4]
  wire [7:0] _T_14697; // @[Mux.scala 46:16:@12161.4]
  wire  _T_14698; // @[Mux.scala 46:19:@12162.4]
  wire [7:0] _T_14699; // @[Mux.scala 46:16:@12163.4]
  wire  _T_14700; // @[Mux.scala 46:19:@12164.4]
  wire [7:0] _T_14701; // @[Mux.scala 46:16:@12165.4]
  wire  _T_14702; // @[Mux.scala 46:19:@12166.4]
  wire [7:0] _T_14703; // @[Mux.scala 46:16:@12167.4]
  wire  _T_14704; // @[Mux.scala 46:19:@12168.4]
  wire [7:0] _T_14705; // @[Mux.scala 46:16:@12169.4]
  wire  _T_14706; // @[Mux.scala 46:19:@12170.4]
  wire [7:0] _T_14707; // @[Mux.scala 46:16:@12171.4]
  wire  _T_14708; // @[Mux.scala 46:19:@12172.4]
  wire [7:0] _T_14709; // @[Mux.scala 46:16:@12173.4]
  wire  _T_14710; // @[Mux.scala 46:19:@12174.4]
  wire [7:0] _T_14711; // @[Mux.scala 46:16:@12175.4]
  wire  _T_14712; // @[Mux.scala 46:19:@12176.4]
  wire [7:0] _T_14713; // @[Mux.scala 46:16:@12177.4]
  wire  _T_14714; // @[Mux.scala 46:19:@12178.4]
  wire [7:0] _T_14715; // @[Mux.scala 46:16:@12179.4]
  wire  _T_14716; // @[Mux.scala 46:19:@12180.4]
  wire [7:0] _T_14717; // @[Mux.scala 46:16:@12181.4]
  wire  _T_14718; // @[Mux.scala 46:19:@12182.4]
  wire [7:0] _T_14719; // @[Mux.scala 46:16:@12183.4]
  wire  _T_14720; // @[Mux.scala 46:19:@12184.4]
  wire [7:0] _T_14721; // @[Mux.scala 46:16:@12185.4]
  wire  _T_14722; // @[Mux.scala 46:19:@12186.4]
  wire [7:0] _T_14723; // @[Mux.scala 46:16:@12187.4]
  wire  _T_14724; // @[Mux.scala 46:19:@12188.4]
  wire [7:0] _T_14725; // @[Mux.scala 46:16:@12189.4]
  wire  _T_14726; // @[Mux.scala 46:19:@12190.4]
  wire [7:0] _T_14727; // @[Mux.scala 46:16:@12191.4]
  wire  _T_14728; // @[Mux.scala 46:19:@12192.4]
  wire [7:0] _T_14729; // @[Mux.scala 46:16:@12193.4]
  wire  _T_14730; // @[Mux.scala 46:19:@12194.4]
  wire [7:0] _T_14731; // @[Mux.scala 46:16:@12195.4]
  wire  _T_14732; // @[Mux.scala 46:19:@12196.4]
  wire [7:0] _T_14733; // @[Mux.scala 46:16:@12197.4]
  wire  _T_14734; // @[Mux.scala 46:19:@12198.4]
  wire [7:0] _T_14735; // @[Mux.scala 46:16:@12199.4]
  wire  _T_14736; // @[Mux.scala 46:19:@12200.4]
  wire [7:0] _T_14737; // @[Mux.scala 46:16:@12201.4]
  wire  _T_14738; // @[Mux.scala 46:19:@12202.4]
  wire [7:0] _T_14739; // @[Mux.scala 46:16:@12203.4]
  wire  _T_14740; // @[Mux.scala 46:19:@12204.4]
  wire [7:0] _T_14741; // @[Mux.scala 46:16:@12205.4]
  wire  _T_14742; // @[Mux.scala 46:19:@12206.4]
  wire [7:0] _T_14743; // @[Mux.scala 46:16:@12207.4]
  wire  _T_14744; // @[Mux.scala 46:19:@12208.4]
  wire [7:0] _T_14745; // @[Mux.scala 46:16:@12209.4]
  wire  _T_14746; // @[Mux.scala 46:19:@12210.4]
  wire [7:0] _T_14747; // @[Mux.scala 46:16:@12211.4]
  wire  _T_14748; // @[Mux.scala 46:19:@12212.4]
  wire [7:0] _T_14749; // @[Mux.scala 46:16:@12213.4]
  wire  _T_14750; // @[Mux.scala 46:19:@12214.4]
  wire [7:0] _T_14751; // @[Mux.scala 46:16:@12215.4]
  wire  _T_14752; // @[Mux.scala 46:19:@12216.4]
  wire [7:0] _T_14753; // @[Mux.scala 46:16:@12217.4]
  wire  _T_14754; // @[Mux.scala 46:19:@12218.4]
  wire [7:0] _T_14755; // @[Mux.scala 46:16:@12219.4]
  wire  _T_14811; // @[Mux.scala 46:19:@12221.4]
  wire [7:0] _T_14812; // @[Mux.scala 46:16:@12222.4]
  wire  _T_14813; // @[Mux.scala 46:19:@12223.4]
  wire [7:0] _T_14814; // @[Mux.scala 46:16:@12224.4]
  wire  _T_14815; // @[Mux.scala 46:19:@12225.4]
  wire [7:0] _T_14816; // @[Mux.scala 46:16:@12226.4]
  wire  _T_14817; // @[Mux.scala 46:19:@12227.4]
  wire [7:0] _T_14818; // @[Mux.scala 46:16:@12228.4]
  wire  _T_14819; // @[Mux.scala 46:19:@12229.4]
  wire [7:0] _T_14820; // @[Mux.scala 46:16:@12230.4]
  wire  _T_14821; // @[Mux.scala 46:19:@12231.4]
  wire [7:0] _T_14822; // @[Mux.scala 46:16:@12232.4]
  wire  _T_14823; // @[Mux.scala 46:19:@12233.4]
  wire [7:0] _T_14824; // @[Mux.scala 46:16:@12234.4]
  wire  _T_14825; // @[Mux.scala 46:19:@12235.4]
  wire [7:0] _T_14826; // @[Mux.scala 46:16:@12236.4]
  wire  _T_14827; // @[Mux.scala 46:19:@12237.4]
  wire [7:0] _T_14828; // @[Mux.scala 46:16:@12238.4]
  wire  _T_14829; // @[Mux.scala 46:19:@12239.4]
  wire [7:0] _T_14830; // @[Mux.scala 46:16:@12240.4]
  wire  _T_14831; // @[Mux.scala 46:19:@12241.4]
  wire [7:0] _T_14832; // @[Mux.scala 46:16:@12242.4]
  wire  _T_14833; // @[Mux.scala 46:19:@12243.4]
  wire [7:0] _T_14834; // @[Mux.scala 46:16:@12244.4]
  wire  _T_14835; // @[Mux.scala 46:19:@12245.4]
  wire [7:0] _T_14836; // @[Mux.scala 46:16:@12246.4]
  wire  _T_14837; // @[Mux.scala 46:19:@12247.4]
  wire [7:0] _T_14838; // @[Mux.scala 46:16:@12248.4]
  wire  _T_14839; // @[Mux.scala 46:19:@12249.4]
  wire [7:0] _T_14840; // @[Mux.scala 46:16:@12250.4]
  wire  _T_14841; // @[Mux.scala 46:19:@12251.4]
  wire [7:0] _T_14842; // @[Mux.scala 46:16:@12252.4]
  wire  _T_14843; // @[Mux.scala 46:19:@12253.4]
  wire [7:0] _T_14844; // @[Mux.scala 46:16:@12254.4]
  wire  _T_14845; // @[Mux.scala 46:19:@12255.4]
  wire [7:0] _T_14846; // @[Mux.scala 46:16:@12256.4]
  wire  _T_14847; // @[Mux.scala 46:19:@12257.4]
  wire [7:0] _T_14848; // @[Mux.scala 46:16:@12258.4]
  wire  _T_14849; // @[Mux.scala 46:19:@12259.4]
  wire [7:0] _T_14850; // @[Mux.scala 46:16:@12260.4]
  wire  _T_14851; // @[Mux.scala 46:19:@12261.4]
  wire [7:0] _T_14852; // @[Mux.scala 46:16:@12262.4]
  wire  _T_14853; // @[Mux.scala 46:19:@12263.4]
  wire [7:0] _T_14854; // @[Mux.scala 46:16:@12264.4]
  wire  _T_14855; // @[Mux.scala 46:19:@12265.4]
  wire [7:0] _T_14856; // @[Mux.scala 46:16:@12266.4]
  wire  _T_14857; // @[Mux.scala 46:19:@12267.4]
  wire [7:0] _T_14858; // @[Mux.scala 46:16:@12268.4]
  wire  _T_14859; // @[Mux.scala 46:19:@12269.4]
  wire [7:0] _T_14860; // @[Mux.scala 46:16:@12270.4]
  wire  _T_14861; // @[Mux.scala 46:19:@12271.4]
  wire [7:0] _T_14862; // @[Mux.scala 46:16:@12272.4]
  wire  _T_14863; // @[Mux.scala 46:19:@12273.4]
  wire [7:0] _T_14864; // @[Mux.scala 46:16:@12274.4]
  wire  _T_14865; // @[Mux.scala 46:19:@12275.4]
  wire [7:0] _T_14866; // @[Mux.scala 46:16:@12276.4]
  wire  _T_14867; // @[Mux.scala 46:19:@12277.4]
  wire [7:0] _T_14868; // @[Mux.scala 46:16:@12278.4]
  wire  _T_14869; // @[Mux.scala 46:19:@12279.4]
  wire [7:0] _T_14870; // @[Mux.scala 46:16:@12280.4]
  wire  _T_14871; // @[Mux.scala 46:19:@12281.4]
  wire [7:0] _T_14872; // @[Mux.scala 46:16:@12282.4]
  wire  _T_14873; // @[Mux.scala 46:19:@12283.4]
  wire [7:0] _T_14874; // @[Mux.scala 46:16:@12284.4]
  wire  _T_14875; // @[Mux.scala 46:19:@12285.4]
  wire [7:0] _T_14876; // @[Mux.scala 46:16:@12286.4]
  wire  _T_14877; // @[Mux.scala 46:19:@12287.4]
  wire [7:0] _T_14878; // @[Mux.scala 46:16:@12288.4]
  wire  _T_14879; // @[Mux.scala 46:19:@12289.4]
  wire [7:0] _T_14880; // @[Mux.scala 46:16:@12290.4]
  wire  _T_14881; // @[Mux.scala 46:19:@12291.4]
  wire [7:0] _T_14882; // @[Mux.scala 46:16:@12292.4]
  wire  _T_14883; // @[Mux.scala 46:19:@12293.4]
  wire [7:0] _T_14884; // @[Mux.scala 46:16:@12294.4]
  wire  _T_14885; // @[Mux.scala 46:19:@12295.4]
  wire [7:0] _T_14886; // @[Mux.scala 46:16:@12296.4]
  wire  _T_14887; // @[Mux.scala 46:19:@12297.4]
  wire [7:0] _T_14888; // @[Mux.scala 46:16:@12298.4]
  wire  _T_14889; // @[Mux.scala 46:19:@12299.4]
  wire [7:0] _T_14890; // @[Mux.scala 46:16:@12300.4]
  wire  _T_14891; // @[Mux.scala 46:19:@12301.4]
  wire [7:0] _T_14892; // @[Mux.scala 46:16:@12302.4]
  wire  _T_14893; // @[Mux.scala 46:19:@12303.4]
  wire [7:0] _T_14894; // @[Mux.scala 46:16:@12304.4]
  wire  _T_14895; // @[Mux.scala 46:19:@12305.4]
  wire [7:0] _T_14896; // @[Mux.scala 46:16:@12306.4]
  wire  _T_14897; // @[Mux.scala 46:19:@12307.4]
  wire [7:0] _T_14898; // @[Mux.scala 46:16:@12308.4]
  wire  _T_14899; // @[Mux.scala 46:19:@12309.4]
  wire [7:0] _T_14900; // @[Mux.scala 46:16:@12310.4]
  wire  _T_14901; // @[Mux.scala 46:19:@12311.4]
  wire [7:0] _T_14902; // @[Mux.scala 46:16:@12312.4]
  wire  _T_14903; // @[Mux.scala 46:19:@12313.4]
  wire [7:0] _T_14904; // @[Mux.scala 46:16:@12314.4]
  wire  _T_14905; // @[Mux.scala 46:19:@12315.4]
  wire [7:0] _T_14906; // @[Mux.scala 46:16:@12316.4]
  wire  _T_14907; // @[Mux.scala 46:19:@12317.4]
  wire [7:0] _T_14908; // @[Mux.scala 46:16:@12318.4]
  wire  _T_14909; // @[Mux.scala 46:19:@12319.4]
  wire [7:0] _T_14910; // @[Mux.scala 46:16:@12320.4]
  wire  _T_14911; // @[Mux.scala 46:19:@12321.4]
  wire [7:0] _T_14912; // @[Mux.scala 46:16:@12322.4]
  wire  _T_14913; // @[Mux.scala 46:19:@12323.4]
  wire [7:0] _T_14914; // @[Mux.scala 46:16:@12324.4]
  wire  _T_14915; // @[Mux.scala 46:19:@12325.4]
  wire [7:0] _T_14916; // @[Mux.scala 46:16:@12326.4]
  wire  _T_14917; // @[Mux.scala 46:19:@12327.4]
  wire [7:0] _T_14918; // @[Mux.scala 46:16:@12328.4]
  wire  _T_14975; // @[Mux.scala 46:19:@12330.4]
  wire [7:0] _T_14976; // @[Mux.scala 46:16:@12331.4]
  wire  _T_14977; // @[Mux.scala 46:19:@12332.4]
  wire [7:0] _T_14978; // @[Mux.scala 46:16:@12333.4]
  wire  _T_14979; // @[Mux.scala 46:19:@12334.4]
  wire [7:0] _T_14980; // @[Mux.scala 46:16:@12335.4]
  wire  _T_14981; // @[Mux.scala 46:19:@12336.4]
  wire [7:0] _T_14982; // @[Mux.scala 46:16:@12337.4]
  wire  _T_14983; // @[Mux.scala 46:19:@12338.4]
  wire [7:0] _T_14984; // @[Mux.scala 46:16:@12339.4]
  wire  _T_14985; // @[Mux.scala 46:19:@12340.4]
  wire [7:0] _T_14986; // @[Mux.scala 46:16:@12341.4]
  wire  _T_14987; // @[Mux.scala 46:19:@12342.4]
  wire [7:0] _T_14988; // @[Mux.scala 46:16:@12343.4]
  wire  _T_14989; // @[Mux.scala 46:19:@12344.4]
  wire [7:0] _T_14990; // @[Mux.scala 46:16:@12345.4]
  wire  _T_14991; // @[Mux.scala 46:19:@12346.4]
  wire [7:0] _T_14992; // @[Mux.scala 46:16:@12347.4]
  wire  _T_14993; // @[Mux.scala 46:19:@12348.4]
  wire [7:0] _T_14994; // @[Mux.scala 46:16:@12349.4]
  wire  _T_14995; // @[Mux.scala 46:19:@12350.4]
  wire [7:0] _T_14996; // @[Mux.scala 46:16:@12351.4]
  wire  _T_14997; // @[Mux.scala 46:19:@12352.4]
  wire [7:0] _T_14998; // @[Mux.scala 46:16:@12353.4]
  wire  _T_14999; // @[Mux.scala 46:19:@12354.4]
  wire [7:0] _T_15000; // @[Mux.scala 46:16:@12355.4]
  wire  _T_15001; // @[Mux.scala 46:19:@12356.4]
  wire [7:0] _T_15002; // @[Mux.scala 46:16:@12357.4]
  wire  _T_15003; // @[Mux.scala 46:19:@12358.4]
  wire [7:0] _T_15004; // @[Mux.scala 46:16:@12359.4]
  wire  _T_15005; // @[Mux.scala 46:19:@12360.4]
  wire [7:0] _T_15006; // @[Mux.scala 46:16:@12361.4]
  wire  _T_15007; // @[Mux.scala 46:19:@12362.4]
  wire [7:0] _T_15008; // @[Mux.scala 46:16:@12363.4]
  wire  _T_15009; // @[Mux.scala 46:19:@12364.4]
  wire [7:0] _T_15010; // @[Mux.scala 46:16:@12365.4]
  wire  _T_15011; // @[Mux.scala 46:19:@12366.4]
  wire [7:0] _T_15012; // @[Mux.scala 46:16:@12367.4]
  wire  _T_15013; // @[Mux.scala 46:19:@12368.4]
  wire [7:0] _T_15014; // @[Mux.scala 46:16:@12369.4]
  wire  _T_15015; // @[Mux.scala 46:19:@12370.4]
  wire [7:0] _T_15016; // @[Mux.scala 46:16:@12371.4]
  wire  _T_15017; // @[Mux.scala 46:19:@12372.4]
  wire [7:0] _T_15018; // @[Mux.scala 46:16:@12373.4]
  wire  _T_15019; // @[Mux.scala 46:19:@12374.4]
  wire [7:0] _T_15020; // @[Mux.scala 46:16:@12375.4]
  wire  _T_15021; // @[Mux.scala 46:19:@12376.4]
  wire [7:0] _T_15022; // @[Mux.scala 46:16:@12377.4]
  wire  _T_15023; // @[Mux.scala 46:19:@12378.4]
  wire [7:0] _T_15024; // @[Mux.scala 46:16:@12379.4]
  wire  _T_15025; // @[Mux.scala 46:19:@12380.4]
  wire [7:0] _T_15026; // @[Mux.scala 46:16:@12381.4]
  wire  _T_15027; // @[Mux.scala 46:19:@12382.4]
  wire [7:0] _T_15028; // @[Mux.scala 46:16:@12383.4]
  wire  _T_15029; // @[Mux.scala 46:19:@12384.4]
  wire [7:0] _T_15030; // @[Mux.scala 46:16:@12385.4]
  wire  _T_15031; // @[Mux.scala 46:19:@12386.4]
  wire [7:0] _T_15032; // @[Mux.scala 46:16:@12387.4]
  wire  _T_15033; // @[Mux.scala 46:19:@12388.4]
  wire [7:0] _T_15034; // @[Mux.scala 46:16:@12389.4]
  wire  _T_15035; // @[Mux.scala 46:19:@12390.4]
  wire [7:0] _T_15036; // @[Mux.scala 46:16:@12391.4]
  wire  _T_15037; // @[Mux.scala 46:19:@12392.4]
  wire [7:0] _T_15038; // @[Mux.scala 46:16:@12393.4]
  wire  _T_15039; // @[Mux.scala 46:19:@12394.4]
  wire [7:0] _T_15040; // @[Mux.scala 46:16:@12395.4]
  wire  _T_15041; // @[Mux.scala 46:19:@12396.4]
  wire [7:0] _T_15042; // @[Mux.scala 46:16:@12397.4]
  wire  _T_15043; // @[Mux.scala 46:19:@12398.4]
  wire [7:0] _T_15044; // @[Mux.scala 46:16:@12399.4]
  wire  _T_15045; // @[Mux.scala 46:19:@12400.4]
  wire [7:0] _T_15046; // @[Mux.scala 46:16:@12401.4]
  wire  _T_15047; // @[Mux.scala 46:19:@12402.4]
  wire [7:0] _T_15048; // @[Mux.scala 46:16:@12403.4]
  wire  _T_15049; // @[Mux.scala 46:19:@12404.4]
  wire [7:0] _T_15050; // @[Mux.scala 46:16:@12405.4]
  wire  _T_15051; // @[Mux.scala 46:19:@12406.4]
  wire [7:0] _T_15052; // @[Mux.scala 46:16:@12407.4]
  wire  _T_15053; // @[Mux.scala 46:19:@12408.4]
  wire [7:0] _T_15054; // @[Mux.scala 46:16:@12409.4]
  wire  _T_15055; // @[Mux.scala 46:19:@12410.4]
  wire [7:0] _T_15056; // @[Mux.scala 46:16:@12411.4]
  wire  _T_15057; // @[Mux.scala 46:19:@12412.4]
  wire [7:0] _T_15058; // @[Mux.scala 46:16:@12413.4]
  wire  _T_15059; // @[Mux.scala 46:19:@12414.4]
  wire [7:0] _T_15060; // @[Mux.scala 46:16:@12415.4]
  wire  _T_15061; // @[Mux.scala 46:19:@12416.4]
  wire [7:0] _T_15062; // @[Mux.scala 46:16:@12417.4]
  wire  _T_15063; // @[Mux.scala 46:19:@12418.4]
  wire [7:0] _T_15064; // @[Mux.scala 46:16:@12419.4]
  wire  _T_15065; // @[Mux.scala 46:19:@12420.4]
  wire [7:0] _T_15066; // @[Mux.scala 46:16:@12421.4]
  wire  _T_15067; // @[Mux.scala 46:19:@12422.4]
  wire [7:0] _T_15068; // @[Mux.scala 46:16:@12423.4]
  wire  _T_15069; // @[Mux.scala 46:19:@12424.4]
  wire [7:0] _T_15070; // @[Mux.scala 46:16:@12425.4]
  wire  _T_15071; // @[Mux.scala 46:19:@12426.4]
  wire [7:0] _T_15072; // @[Mux.scala 46:16:@12427.4]
  wire  _T_15073; // @[Mux.scala 46:19:@12428.4]
  wire [7:0] _T_15074; // @[Mux.scala 46:16:@12429.4]
  wire  _T_15075; // @[Mux.scala 46:19:@12430.4]
  wire [7:0] _T_15076; // @[Mux.scala 46:16:@12431.4]
  wire  _T_15077; // @[Mux.scala 46:19:@12432.4]
  wire [7:0] _T_15078; // @[Mux.scala 46:16:@12433.4]
  wire  _T_15079; // @[Mux.scala 46:19:@12434.4]
  wire [7:0] _T_15080; // @[Mux.scala 46:16:@12435.4]
  wire  _T_15081; // @[Mux.scala 46:19:@12436.4]
  wire [7:0] _T_15082; // @[Mux.scala 46:16:@12437.4]
  wire  _T_15083; // @[Mux.scala 46:19:@12438.4]
  wire [7:0] _T_15084; // @[Mux.scala 46:16:@12439.4]
  wire  _T_15142; // @[Mux.scala 46:19:@12441.4]
  wire [7:0] _T_15143; // @[Mux.scala 46:16:@12442.4]
  wire  _T_15144; // @[Mux.scala 46:19:@12443.4]
  wire [7:0] _T_15145; // @[Mux.scala 46:16:@12444.4]
  wire  _T_15146; // @[Mux.scala 46:19:@12445.4]
  wire [7:0] _T_15147; // @[Mux.scala 46:16:@12446.4]
  wire  _T_15148; // @[Mux.scala 46:19:@12447.4]
  wire [7:0] _T_15149; // @[Mux.scala 46:16:@12448.4]
  wire  _T_15150; // @[Mux.scala 46:19:@12449.4]
  wire [7:0] _T_15151; // @[Mux.scala 46:16:@12450.4]
  wire  _T_15152; // @[Mux.scala 46:19:@12451.4]
  wire [7:0] _T_15153; // @[Mux.scala 46:16:@12452.4]
  wire  _T_15154; // @[Mux.scala 46:19:@12453.4]
  wire [7:0] _T_15155; // @[Mux.scala 46:16:@12454.4]
  wire  _T_15156; // @[Mux.scala 46:19:@12455.4]
  wire [7:0] _T_15157; // @[Mux.scala 46:16:@12456.4]
  wire  _T_15158; // @[Mux.scala 46:19:@12457.4]
  wire [7:0] _T_15159; // @[Mux.scala 46:16:@12458.4]
  wire  _T_15160; // @[Mux.scala 46:19:@12459.4]
  wire [7:0] _T_15161; // @[Mux.scala 46:16:@12460.4]
  wire  _T_15162; // @[Mux.scala 46:19:@12461.4]
  wire [7:0] _T_15163; // @[Mux.scala 46:16:@12462.4]
  wire  _T_15164; // @[Mux.scala 46:19:@12463.4]
  wire [7:0] _T_15165; // @[Mux.scala 46:16:@12464.4]
  wire  _T_15166; // @[Mux.scala 46:19:@12465.4]
  wire [7:0] _T_15167; // @[Mux.scala 46:16:@12466.4]
  wire  _T_15168; // @[Mux.scala 46:19:@12467.4]
  wire [7:0] _T_15169; // @[Mux.scala 46:16:@12468.4]
  wire  _T_15170; // @[Mux.scala 46:19:@12469.4]
  wire [7:0] _T_15171; // @[Mux.scala 46:16:@12470.4]
  wire  _T_15172; // @[Mux.scala 46:19:@12471.4]
  wire [7:0] _T_15173; // @[Mux.scala 46:16:@12472.4]
  wire  _T_15174; // @[Mux.scala 46:19:@12473.4]
  wire [7:0] _T_15175; // @[Mux.scala 46:16:@12474.4]
  wire  _T_15176; // @[Mux.scala 46:19:@12475.4]
  wire [7:0] _T_15177; // @[Mux.scala 46:16:@12476.4]
  wire  _T_15178; // @[Mux.scala 46:19:@12477.4]
  wire [7:0] _T_15179; // @[Mux.scala 46:16:@12478.4]
  wire  _T_15180; // @[Mux.scala 46:19:@12479.4]
  wire [7:0] _T_15181; // @[Mux.scala 46:16:@12480.4]
  wire  _T_15182; // @[Mux.scala 46:19:@12481.4]
  wire [7:0] _T_15183; // @[Mux.scala 46:16:@12482.4]
  wire  _T_15184; // @[Mux.scala 46:19:@12483.4]
  wire [7:0] _T_15185; // @[Mux.scala 46:16:@12484.4]
  wire  _T_15186; // @[Mux.scala 46:19:@12485.4]
  wire [7:0] _T_15187; // @[Mux.scala 46:16:@12486.4]
  wire  _T_15188; // @[Mux.scala 46:19:@12487.4]
  wire [7:0] _T_15189; // @[Mux.scala 46:16:@12488.4]
  wire  _T_15190; // @[Mux.scala 46:19:@12489.4]
  wire [7:0] _T_15191; // @[Mux.scala 46:16:@12490.4]
  wire  _T_15192; // @[Mux.scala 46:19:@12491.4]
  wire [7:0] _T_15193; // @[Mux.scala 46:16:@12492.4]
  wire  _T_15194; // @[Mux.scala 46:19:@12493.4]
  wire [7:0] _T_15195; // @[Mux.scala 46:16:@12494.4]
  wire  _T_15196; // @[Mux.scala 46:19:@12495.4]
  wire [7:0] _T_15197; // @[Mux.scala 46:16:@12496.4]
  wire  _T_15198; // @[Mux.scala 46:19:@12497.4]
  wire [7:0] _T_15199; // @[Mux.scala 46:16:@12498.4]
  wire  _T_15200; // @[Mux.scala 46:19:@12499.4]
  wire [7:0] _T_15201; // @[Mux.scala 46:16:@12500.4]
  wire  _T_15202; // @[Mux.scala 46:19:@12501.4]
  wire [7:0] _T_15203; // @[Mux.scala 46:16:@12502.4]
  wire  _T_15204; // @[Mux.scala 46:19:@12503.4]
  wire [7:0] _T_15205; // @[Mux.scala 46:16:@12504.4]
  wire  _T_15206; // @[Mux.scala 46:19:@12505.4]
  wire [7:0] _T_15207; // @[Mux.scala 46:16:@12506.4]
  wire  _T_15208; // @[Mux.scala 46:19:@12507.4]
  wire [7:0] _T_15209; // @[Mux.scala 46:16:@12508.4]
  wire  _T_15210; // @[Mux.scala 46:19:@12509.4]
  wire [7:0] _T_15211; // @[Mux.scala 46:16:@12510.4]
  wire  _T_15212; // @[Mux.scala 46:19:@12511.4]
  wire [7:0] _T_15213; // @[Mux.scala 46:16:@12512.4]
  wire  _T_15214; // @[Mux.scala 46:19:@12513.4]
  wire [7:0] _T_15215; // @[Mux.scala 46:16:@12514.4]
  wire  _T_15216; // @[Mux.scala 46:19:@12515.4]
  wire [7:0] _T_15217; // @[Mux.scala 46:16:@12516.4]
  wire  _T_15218; // @[Mux.scala 46:19:@12517.4]
  wire [7:0] _T_15219; // @[Mux.scala 46:16:@12518.4]
  wire  _T_15220; // @[Mux.scala 46:19:@12519.4]
  wire [7:0] _T_15221; // @[Mux.scala 46:16:@12520.4]
  wire  _T_15222; // @[Mux.scala 46:19:@12521.4]
  wire [7:0] _T_15223; // @[Mux.scala 46:16:@12522.4]
  wire  _T_15224; // @[Mux.scala 46:19:@12523.4]
  wire [7:0] _T_15225; // @[Mux.scala 46:16:@12524.4]
  wire  _T_15226; // @[Mux.scala 46:19:@12525.4]
  wire [7:0] _T_15227; // @[Mux.scala 46:16:@12526.4]
  wire  _T_15228; // @[Mux.scala 46:19:@12527.4]
  wire [7:0] _T_15229; // @[Mux.scala 46:16:@12528.4]
  wire  _T_15230; // @[Mux.scala 46:19:@12529.4]
  wire [7:0] _T_15231; // @[Mux.scala 46:16:@12530.4]
  wire  _T_15232; // @[Mux.scala 46:19:@12531.4]
  wire [7:0] _T_15233; // @[Mux.scala 46:16:@12532.4]
  wire  _T_15234; // @[Mux.scala 46:19:@12533.4]
  wire [7:0] _T_15235; // @[Mux.scala 46:16:@12534.4]
  wire  _T_15236; // @[Mux.scala 46:19:@12535.4]
  wire [7:0] _T_15237; // @[Mux.scala 46:16:@12536.4]
  wire  _T_15238; // @[Mux.scala 46:19:@12537.4]
  wire [7:0] _T_15239; // @[Mux.scala 46:16:@12538.4]
  wire  _T_15240; // @[Mux.scala 46:19:@12539.4]
  wire [7:0] _T_15241; // @[Mux.scala 46:16:@12540.4]
  wire  _T_15242; // @[Mux.scala 46:19:@12541.4]
  wire [7:0] _T_15243; // @[Mux.scala 46:16:@12542.4]
  wire  _T_15244; // @[Mux.scala 46:19:@12543.4]
  wire [7:0] _T_15245; // @[Mux.scala 46:16:@12544.4]
  wire  _T_15246; // @[Mux.scala 46:19:@12545.4]
  wire [7:0] _T_15247; // @[Mux.scala 46:16:@12546.4]
  wire  _T_15248; // @[Mux.scala 46:19:@12547.4]
  wire [7:0] _T_15249; // @[Mux.scala 46:16:@12548.4]
  wire  _T_15250; // @[Mux.scala 46:19:@12549.4]
  wire [7:0] _T_15251; // @[Mux.scala 46:16:@12550.4]
  wire  _T_15252; // @[Mux.scala 46:19:@12551.4]
  wire [7:0] _T_15253; // @[Mux.scala 46:16:@12552.4]
  wire  _T_15312; // @[Mux.scala 46:19:@12554.4]
  wire [7:0] _T_15313; // @[Mux.scala 46:16:@12555.4]
  wire  _T_15314; // @[Mux.scala 46:19:@12556.4]
  wire [7:0] _T_15315; // @[Mux.scala 46:16:@12557.4]
  wire  _T_15316; // @[Mux.scala 46:19:@12558.4]
  wire [7:0] _T_15317; // @[Mux.scala 46:16:@12559.4]
  wire  _T_15318; // @[Mux.scala 46:19:@12560.4]
  wire [7:0] _T_15319; // @[Mux.scala 46:16:@12561.4]
  wire  _T_15320; // @[Mux.scala 46:19:@12562.4]
  wire [7:0] _T_15321; // @[Mux.scala 46:16:@12563.4]
  wire  _T_15322; // @[Mux.scala 46:19:@12564.4]
  wire [7:0] _T_15323; // @[Mux.scala 46:16:@12565.4]
  wire  _T_15324; // @[Mux.scala 46:19:@12566.4]
  wire [7:0] _T_15325; // @[Mux.scala 46:16:@12567.4]
  wire  _T_15326; // @[Mux.scala 46:19:@12568.4]
  wire [7:0] _T_15327; // @[Mux.scala 46:16:@12569.4]
  wire  _T_15328; // @[Mux.scala 46:19:@12570.4]
  wire [7:0] _T_15329; // @[Mux.scala 46:16:@12571.4]
  wire  _T_15330; // @[Mux.scala 46:19:@12572.4]
  wire [7:0] _T_15331; // @[Mux.scala 46:16:@12573.4]
  wire  _T_15332; // @[Mux.scala 46:19:@12574.4]
  wire [7:0] _T_15333; // @[Mux.scala 46:16:@12575.4]
  wire  _T_15334; // @[Mux.scala 46:19:@12576.4]
  wire [7:0] _T_15335; // @[Mux.scala 46:16:@12577.4]
  wire  _T_15336; // @[Mux.scala 46:19:@12578.4]
  wire [7:0] _T_15337; // @[Mux.scala 46:16:@12579.4]
  wire  _T_15338; // @[Mux.scala 46:19:@12580.4]
  wire [7:0] _T_15339; // @[Mux.scala 46:16:@12581.4]
  wire  _T_15340; // @[Mux.scala 46:19:@12582.4]
  wire [7:0] _T_15341; // @[Mux.scala 46:16:@12583.4]
  wire  _T_15342; // @[Mux.scala 46:19:@12584.4]
  wire [7:0] _T_15343; // @[Mux.scala 46:16:@12585.4]
  wire  _T_15344; // @[Mux.scala 46:19:@12586.4]
  wire [7:0] _T_15345; // @[Mux.scala 46:16:@12587.4]
  wire  _T_15346; // @[Mux.scala 46:19:@12588.4]
  wire [7:0] _T_15347; // @[Mux.scala 46:16:@12589.4]
  wire  _T_15348; // @[Mux.scala 46:19:@12590.4]
  wire [7:0] _T_15349; // @[Mux.scala 46:16:@12591.4]
  wire  _T_15350; // @[Mux.scala 46:19:@12592.4]
  wire [7:0] _T_15351; // @[Mux.scala 46:16:@12593.4]
  wire  _T_15352; // @[Mux.scala 46:19:@12594.4]
  wire [7:0] _T_15353; // @[Mux.scala 46:16:@12595.4]
  wire  _T_15354; // @[Mux.scala 46:19:@12596.4]
  wire [7:0] _T_15355; // @[Mux.scala 46:16:@12597.4]
  wire  _T_15356; // @[Mux.scala 46:19:@12598.4]
  wire [7:0] _T_15357; // @[Mux.scala 46:16:@12599.4]
  wire  _T_15358; // @[Mux.scala 46:19:@12600.4]
  wire [7:0] _T_15359; // @[Mux.scala 46:16:@12601.4]
  wire  _T_15360; // @[Mux.scala 46:19:@12602.4]
  wire [7:0] _T_15361; // @[Mux.scala 46:16:@12603.4]
  wire  _T_15362; // @[Mux.scala 46:19:@12604.4]
  wire [7:0] _T_15363; // @[Mux.scala 46:16:@12605.4]
  wire  _T_15364; // @[Mux.scala 46:19:@12606.4]
  wire [7:0] _T_15365; // @[Mux.scala 46:16:@12607.4]
  wire  _T_15366; // @[Mux.scala 46:19:@12608.4]
  wire [7:0] _T_15367; // @[Mux.scala 46:16:@12609.4]
  wire  _T_15368; // @[Mux.scala 46:19:@12610.4]
  wire [7:0] _T_15369; // @[Mux.scala 46:16:@12611.4]
  wire  _T_15370; // @[Mux.scala 46:19:@12612.4]
  wire [7:0] _T_15371; // @[Mux.scala 46:16:@12613.4]
  wire  _T_15372; // @[Mux.scala 46:19:@12614.4]
  wire [7:0] _T_15373; // @[Mux.scala 46:16:@12615.4]
  wire  _T_15374; // @[Mux.scala 46:19:@12616.4]
  wire [7:0] _T_15375; // @[Mux.scala 46:16:@12617.4]
  wire  _T_15376; // @[Mux.scala 46:19:@12618.4]
  wire [7:0] _T_15377; // @[Mux.scala 46:16:@12619.4]
  wire  _T_15378; // @[Mux.scala 46:19:@12620.4]
  wire [7:0] _T_15379; // @[Mux.scala 46:16:@12621.4]
  wire  _T_15380; // @[Mux.scala 46:19:@12622.4]
  wire [7:0] _T_15381; // @[Mux.scala 46:16:@12623.4]
  wire  _T_15382; // @[Mux.scala 46:19:@12624.4]
  wire [7:0] _T_15383; // @[Mux.scala 46:16:@12625.4]
  wire  _T_15384; // @[Mux.scala 46:19:@12626.4]
  wire [7:0] _T_15385; // @[Mux.scala 46:16:@12627.4]
  wire  _T_15386; // @[Mux.scala 46:19:@12628.4]
  wire [7:0] _T_15387; // @[Mux.scala 46:16:@12629.4]
  wire  _T_15388; // @[Mux.scala 46:19:@12630.4]
  wire [7:0] _T_15389; // @[Mux.scala 46:16:@12631.4]
  wire  _T_15390; // @[Mux.scala 46:19:@12632.4]
  wire [7:0] _T_15391; // @[Mux.scala 46:16:@12633.4]
  wire  _T_15392; // @[Mux.scala 46:19:@12634.4]
  wire [7:0] _T_15393; // @[Mux.scala 46:16:@12635.4]
  wire  _T_15394; // @[Mux.scala 46:19:@12636.4]
  wire [7:0] _T_15395; // @[Mux.scala 46:16:@12637.4]
  wire  _T_15396; // @[Mux.scala 46:19:@12638.4]
  wire [7:0] _T_15397; // @[Mux.scala 46:16:@12639.4]
  wire  _T_15398; // @[Mux.scala 46:19:@12640.4]
  wire [7:0] _T_15399; // @[Mux.scala 46:16:@12641.4]
  wire  _T_15400; // @[Mux.scala 46:19:@12642.4]
  wire [7:0] _T_15401; // @[Mux.scala 46:16:@12643.4]
  wire  _T_15402; // @[Mux.scala 46:19:@12644.4]
  wire [7:0] _T_15403; // @[Mux.scala 46:16:@12645.4]
  wire  _T_15404; // @[Mux.scala 46:19:@12646.4]
  wire [7:0] _T_15405; // @[Mux.scala 46:16:@12647.4]
  wire  _T_15406; // @[Mux.scala 46:19:@12648.4]
  wire [7:0] _T_15407; // @[Mux.scala 46:16:@12649.4]
  wire  _T_15408; // @[Mux.scala 46:19:@12650.4]
  wire [7:0] _T_15409; // @[Mux.scala 46:16:@12651.4]
  wire  _T_15410; // @[Mux.scala 46:19:@12652.4]
  wire [7:0] _T_15411; // @[Mux.scala 46:16:@12653.4]
  wire  _T_15412; // @[Mux.scala 46:19:@12654.4]
  wire [7:0] _T_15413; // @[Mux.scala 46:16:@12655.4]
  wire  _T_15414; // @[Mux.scala 46:19:@12656.4]
  wire [7:0] _T_15415; // @[Mux.scala 46:16:@12657.4]
  wire  _T_15416; // @[Mux.scala 46:19:@12658.4]
  wire [7:0] _T_15417; // @[Mux.scala 46:16:@12659.4]
  wire  _T_15418; // @[Mux.scala 46:19:@12660.4]
  wire [7:0] _T_15419; // @[Mux.scala 46:16:@12661.4]
  wire  _T_15420; // @[Mux.scala 46:19:@12662.4]
  wire [7:0] _T_15421; // @[Mux.scala 46:16:@12663.4]
  wire  _T_15422; // @[Mux.scala 46:19:@12664.4]
  wire [7:0] _T_15423; // @[Mux.scala 46:16:@12665.4]
  wire  _T_15424; // @[Mux.scala 46:19:@12666.4]
  wire [7:0] _T_15425; // @[Mux.scala 46:16:@12667.4]
  wire  _T_15485; // @[Mux.scala 46:19:@12669.4]
  wire [7:0] _T_15486; // @[Mux.scala 46:16:@12670.4]
  wire  _T_15487; // @[Mux.scala 46:19:@12671.4]
  wire [7:0] _T_15488; // @[Mux.scala 46:16:@12672.4]
  wire  _T_15489; // @[Mux.scala 46:19:@12673.4]
  wire [7:0] _T_15490; // @[Mux.scala 46:16:@12674.4]
  wire  _T_15491; // @[Mux.scala 46:19:@12675.4]
  wire [7:0] _T_15492; // @[Mux.scala 46:16:@12676.4]
  wire  _T_15493; // @[Mux.scala 46:19:@12677.4]
  wire [7:0] _T_15494; // @[Mux.scala 46:16:@12678.4]
  wire  _T_15495; // @[Mux.scala 46:19:@12679.4]
  wire [7:0] _T_15496; // @[Mux.scala 46:16:@12680.4]
  wire  _T_15497; // @[Mux.scala 46:19:@12681.4]
  wire [7:0] _T_15498; // @[Mux.scala 46:16:@12682.4]
  wire  _T_15499; // @[Mux.scala 46:19:@12683.4]
  wire [7:0] _T_15500; // @[Mux.scala 46:16:@12684.4]
  wire  _T_15501; // @[Mux.scala 46:19:@12685.4]
  wire [7:0] _T_15502; // @[Mux.scala 46:16:@12686.4]
  wire  _T_15503; // @[Mux.scala 46:19:@12687.4]
  wire [7:0] _T_15504; // @[Mux.scala 46:16:@12688.4]
  wire  _T_15505; // @[Mux.scala 46:19:@12689.4]
  wire [7:0] _T_15506; // @[Mux.scala 46:16:@12690.4]
  wire  _T_15507; // @[Mux.scala 46:19:@12691.4]
  wire [7:0] _T_15508; // @[Mux.scala 46:16:@12692.4]
  wire  _T_15509; // @[Mux.scala 46:19:@12693.4]
  wire [7:0] _T_15510; // @[Mux.scala 46:16:@12694.4]
  wire  _T_15511; // @[Mux.scala 46:19:@12695.4]
  wire [7:0] _T_15512; // @[Mux.scala 46:16:@12696.4]
  wire  _T_15513; // @[Mux.scala 46:19:@12697.4]
  wire [7:0] _T_15514; // @[Mux.scala 46:16:@12698.4]
  wire  _T_15515; // @[Mux.scala 46:19:@12699.4]
  wire [7:0] _T_15516; // @[Mux.scala 46:16:@12700.4]
  wire  _T_15517; // @[Mux.scala 46:19:@12701.4]
  wire [7:0] _T_15518; // @[Mux.scala 46:16:@12702.4]
  wire  _T_15519; // @[Mux.scala 46:19:@12703.4]
  wire [7:0] _T_15520; // @[Mux.scala 46:16:@12704.4]
  wire  _T_15521; // @[Mux.scala 46:19:@12705.4]
  wire [7:0] _T_15522; // @[Mux.scala 46:16:@12706.4]
  wire  _T_15523; // @[Mux.scala 46:19:@12707.4]
  wire [7:0] _T_15524; // @[Mux.scala 46:16:@12708.4]
  wire  _T_15525; // @[Mux.scala 46:19:@12709.4]
  wire [7:0] _T_15526; // @[Mux.scala 46:16:@12710.4]
  wire  _T_15527; // @[Mux.scala 46:19:@12711.4]
  wire [7:0] _T_15528; // @[Mux.scala 46:16:@12712.4]
  wire  _T_15529; // @[Mux.scala 46:19:@12713.4]
  wire [7:0] _T_15530; // @[Mux.scala 46:16:@12714.4]
  wire  _T_15531; // @[Mux.scala 46:19:@12715.4]
  wire [7:0] _T_15532; // @[Mux.scala 46:16:@12716.4]
  wire  _T_15533; // @[Mux.scala 46:19:@12717.4]
  wire [7:0] _T_15534; // @[Mux.scala 46:16:@12718.4]
  wire  _T_15535; // @[Mux.scala 46:19:@12719.4]
  wire [7:0] _T_15536; // @[Mux.scala 46:16:@12720.4]
  wire  _T_15537; // @[Mux.scala 46:19:@12721.4]
  wire [7:0] _T_15538; // @[Mux.scala 46:16:@12722.4]
  wire  _T_15539; // @[Mux.scala 46:19:@12723.4]
  wire [7:0] _T_15540; // @[Mux.scala 46:16:@12724.4]
  wire  _T_15541; // @[Mux.scala 46:19:@12725.4]
  wire [7:0] _T_15542; // @[Mux.scala 46:16:@12726.4]
  wire  _T_15543; // @[Mux.scala 46:19:@12727.4]
  wire [7:0] _T_15544; // @[Mux.scala 46:16:@12728.4]
  wire  _T_15545; // @[Mux.scala 46:19:@12729.4]
  wire [7:0] _T_15546; // @[Mux.scala 46:16:@12730.4]
  wire  _T_15547; // @[Mux.scala 46:19:@12731.4]
  wire [7:0] _T_15548; // @[Mux.scala 46:16:@12732.4]
  wire  _T_15549; // @[Mux.scala 46:19:@12733.4]
  wire [7:0] _T_15550; // @[Mux.scala 46:16:@12734.4]
  wire  _T_15551; // @[Mux.scala 46:19:@12735.4]
  wire [7:0] _T_15552; // @[Mux.scala 46:16:@12736.4]
  wire  _T_15553; // @[Mux.scala 46:19:@12737.4]
  wire [7:0] _T_15554; // @[Mux.scala 46:16:@12738.4]
  wire  _T_15555; // @[Mux.scala 46:19:@12739.4]
  wire [7:0] _T_15556; // @[Mux.scala 46:16:@12740.4]
  wire  _T_15557; // @[Mux.scala 46:19:@12741.4]
  wire [7:0] _T_15558; // @[Mux.scala 46:16:@12742.4]
  wire  _T_15559; // @[Mux.scala 46:19:@12743.4]
  wire [7:0] _T_15560; // @[Mux.scala 46:16:@12744.4]
  wire  _T_15561; // @[Mux.scala 46:19:@12745.4]
  wire [7:0] _T_15562; // @[Mux.scala 46:16:@12746.4]
  wire  _T_15563; // @[Mux.scala 46:19:@12747.4]
  wire [7:0] _T_15564; // @[Mux.scala 46:16:@12748.4]
  wire  _T_15565; // @[Mux.scala 46:19:@12749.4]
  wire [7:0] _T_15566; // @[Mux.scala 46:16:@12750.4]
  wire  _T_15567; // @[Mux.scala 46:19:@12751.4]
  wire [7:0] _T_15568; // @[Mux.scala 46:16:@12752.4]
  wire  _T_15569; // @[Mux.scala 46:19:@12753.4]
  wire [7:0] _T_15570; // @[Mux.scala 46:16:@12754.4]
  wire  _T_15571; // @[Mux.scala 46:19:@12755.4]
  wire [7:0] _T_15572; // @[Mux.scala 46:16:@12756.4]
  wire  _T_15573; // @[Mux.scala 46:19:@12757.4]
  wire [7:0] _T_15574; // @[Mux.scala 46:16:@12758.4]
  wire  _T_15575; // @[Mux.scala 46:19:@12759.4]
  wire [7:0] _T_15576; // @[Mux.scala 46:16:@12760.4]
  wire  _T_15577; // @[Mux.scala 46:19:@12761.4]
  wire [7:0] _T_15578; // @[Mux.scala 46:16:@12762.4]
  wire  _T_15579; // @[Mux.scala 46:19:@12763.4]
  wire [7:0] _T_15580; // @[Mux.scala 46:16:@12764.4]
  wire  _T_15581; // @[Mux.scala 46:19:@12765.4]
  wire [7:0] _T_15582; // @[Mux.scala 46:16:@12766.4]
  wire  _T_15583; // @[Mux.scala 46:19:@12767.4]
  wire [7:0] _T_15584; // @[Mux.scala 46:16:@12768.4]
  wire  _T_15585; // @[Mux.scala 46:19:@12769.4]
  wire [7:0] _T_15586; // @[Mux.scala 46:16:@12770.4]
  wire  _T_15587; // @[Mux.scala 46:19:@12771.4]
  wire [7:0] _T_15588; // @[Mux.scala 46:16:@12772.4]
  wire  _T_15589; // @[Mux.scala 46:19:@12773.4]
  wire [7:0] _T_15590; // @[Mux.scala 46:16:@12774.4]
  wire  _T_15591; // @[Mux.scala 46:19:@12775.4]
  wire [7:0] _T_15592; // @[Mux.scala 46:16:@12776.4]
  wire  _T_15593; // @[Mux.scala 46:19:@12777.4]
  wire [7:0] _T_15594; // @[Mux.scala 46:16:@12778.4]
  wire  _T_15595; // @[Mux.scala 46:19:@12779.4]
  wire [7:0] _T_15596; // @[Mux.scala 46:16:@12780.4]
  wire  _T_15597; // @[Mux.scala 46:19:@12781.4]
  wire [7:0] _T_15598; // @[Mux.scala 46:16:@12782.4]
  wire  _T_15599; // @[Mux.scala 46:19:@12783.4]
  wire [7:0] _T_15600; // @[Mux.scala 46:16:@12784.4]
  wire  _T_15661; // @[Mux.scala 46:19:@12786.4]
  wire [7:0] _T_15662; // @[Mux.scala 46:16:@12787.4]
  wire  _T_15663; // @[Mux.scala 46:19:@12788.4]
  wire [7:0] _T_15664; // @[Mux.scala 46:16:@12789.4]
  wire  _T_15665; // @[Mux.scala 46:19:@12790.4]
  wire [7:0] _T_15666; // @[Mux.scala 46:16:@12791.4]
  wire  _T_15667; // @[Mux.scala 46:19:@12792.4]
  wire [7:0] _T_15668; // @[Mux.scala 46:16:@12793.4]
  wire  _T_15669; // @[Mux.scala 46:19:@12794.4]
  wire [7:0] _T_15670; // @[Mux.scala 46:16:@12795.4]
  wire  _T_15671; // @[Mux.scala 46:19:@12796.4]
  wire [7:0] _T_15672; // @[Mux.scala 46:16:@12797.4]
  wire  _T_15673; // @[Mux.scala 46:19:@12798.4]
  wire [7:0] _T_15674; // @[Mux.scala 46:16:@12799.4]
  wire  _T_15675; // @[Mux.scala 46:19:@12800.4]
  wire [7:0] _T_15676; // @[Mux.scala 46:16:@12801.4]
  wire  _T_15677; // @[Mux.scala 46:19:@12802.4]
  wire [7:0] _T_15678; // @[Mux.scala 46:16:@12803.4]
  wire  _T_15679; // @[Mux.scala 46:19:@12804.4]
  wire [7:0] _T_15680; // @[Mux.scala 46:16:@12805.4]
  wire  _T_15681; // @[Mux.scala 46:19:@12806.4]
  wire [7:0] _T_15682; // @[Mux.scala 46:16:@12807.4]
  wire  _T_15683; // @[Mux.scala 46:19:@12808.4]
  wire [7:0] _T_15684; // @[Mux.scala 46:16:@12809.4]
  wire  _T_15685; // @[Mux.scala 46:19:@12810.4]
  wire [7:0] _T_15686; // @[Mux.scala 46:16:@12811.4]
  wire  _T_15687; // @[Mux.scala 46:19:@12812.4]
  wire [7:0] _T_15688; // @[Mux.scala 46:16:@12813.4]
  wire  _T_15689; // @[Mux.scala 46:19:@12814.4]
  wire [7:0] _T_15690; // @[Mux.scala 46:16:@12815.4]
  wire  _T_15691; // @[Mux.scala 46:19:@12816.4]
  wire [7:0] _T_15692; // @[Mux.scala 46:16:@12817.4]
  wire  _T_15693; // @[Mux.scala 46:19:@12818.4]
  wire [7:0] _T_15694; // @[Mux.scala 46:16:@12819.4]
  wire  _T_15695; // @[Mux.scala 46:19:@12820.4]
  wire [7:0] _T_15696; // @[Mux.scala 46:16:@12821.4]
  wire  _T_15697; // @[Mux.scala 46:19:@12822.4]
  wire [7:0] _T_15698; // @[Mux.scala 46:16:@12823.4]
  wire  _T_15699; // @[Mux.scala 46:19:@12824.4]
  wire [7:0] _T_15700; // @[Mux.scala 46:16:@12825.4]
  wire  _T_15701; // @[Mux.scala 46:19:@12826.4]
  wire [7:0] _T_15702; // @[Mux.scala 46:16:@12827.4]
  wire  _T_15703; // @[Mux.scala 46:19:@12828.4]
  wire [7:0] _T_15704; // @[Mux.scala 46:16:@12829.4]
  wire  _T_15705; // @[Mux.scala 46:19:@12830.4]
  wire [7:0] _T_15706; // @[Mux.scala 46:16:@12831.4]
  wire  _T_15707; // @[Mux.scala 46:19:@12832.4]
  wire [7:0] _T_15708; // @[Mux.scala 46:16:@12833.4]
  wire  _T_15709; // @[Mux.scala 46:19:@12834.4]
  wire [7:0] _T_15710; // @[Mux.scala 46:16:@12835.4]
  wire  _T_15711; // @[Mux.scala 46:19:@12836.4]
  wire [7:0] _T_15712; // @[Mux.scala 46:16:@12837.4]
  wire  _T_15713; // @[Mux.scala 46:19:@12838.4]
  wire [7:0] _T_15714; // @[Mux.scala 46:16:@12839.4]
  wire  _T_15715; // @[Mux.scala 46:19:@12840.4]
  wire [7:0] _T_15716; // @[Mux.scala 46:16:@12841.4]
  wire  _T_15717; // @[Mux.scala 46:19:@12842.4]
  wire [7:0] _T_15718; // @[Mux.scala 46:16:@12843.4]
  wire  _T_15719; // @[Mux.scala 46:19:@12844.4]
  wire [7:0] _T_15720; // @[Mux.scala 46:16:@12845.4]
  wire  _T_15721; // @[Mux.scala 46:19:@12846.4]
  wire [7:0] _T_15722; // @[Mux.scala 46:16:@12847.4]
  wire  _T_15723; // @[Mux.scala 46:19:@12848.4]
  wire [7:0] _T_15724; // @[Mux.scala 46:16:@12849.4]
  wire  _T_15725; // @[Mux.scala 46:19:@12850.4]
  wire [7:0] _T_15726; // @[Mux.scala 46:16:@12851.4]
  wire  _T_15727; // @[Mux.scala 46:19:@12852.4]
  wire [7:0] _T_15728; // @[Mux.scala 46:16:@12853.4]
  wire  _T_15729; // @[Mux.scala 46:19:@12854.4]
  wire [7:0] _T_15730; // @[Mux.scala 46:16:@12855.4]
  wire  _T_15731; // @[Mux.scala 46:19:@12856.4]
  wire [7:0] _T_15732; // @[Mux.scala 46:16:@12857.4]
  wire  _T_15733; // @[Mux.scala 46:19:@12858.4]
  wire [7:0] _T_15734; // @[Mux.scala 46:16:@12859.4]
  wire  _T_15735; // @[Mux.scala 46:19:@12860.4]
  wire [7:0] _T_15736; // @[Mux.scala 46:16:@12861.4]
  wire  _T_15737; // @[Mux.scala 46:19:@12862.4]
  wire [7:0] _T_15738; // @[Mux.scala 46:16:@12863.4]
  wire  _T_15739; // @[Mux.scala 46:19:@12864.4]
  wire [7:0] _T_15740; // @[Mux.scala 46:16:@12865.4]
  wire  _T_15741; // @[Mux.scala 46:19:@12866.4]
  wire [7:0] _T_15742; // @[Mux.scala 46:16:@12867.4]
  wire  _T_15743; // @[Mux.scala 46:19:@12868.4]
  wire [7:0] _T_15744; // @[Mux.scala 46:16:@12869.4]
  wire  _T_15745; // @[Mux.scala 46:19:@12870.4]
  wire [7:0] _T_15746; // @[Mux.scala 46:16:@12871.4]
  wire  _T_15747; // @[Mux.scala 46:19:@12872.4]
  wire [7:0] _T_15748; // @[Mux.scala 46:16:@12873.4]
  wire  _T_15749; // @[Mux.scala 46:19:@12874.4]
  wire [7:0] _T_15750; // @[Mux.scala 46:16:@12875.4]
  wire  _T_15751; // @[Mux.scala 46:19:@12876.4]
  wire [7:0] _T_15752; // @[Mux.scala 46:16:@12877.4]
  wire  _T_15753; // @[Mux.scala 46:19:@12878.4]
  wire [7:0] _T_15754; // @[Mux.scala 46:16:@12879.4]
  wire  _T_15755; // @[Mux.scala 46:19:@12880.4]
  wire [7:0] _T_15756; // @[Mux.scala 46:16:@12881.4]
  wire  _T_15757; // @[Mux.scala 46:19:@12882.4]
  wire [7:0] _T_15758; // @[Mux.scala 46:16:@12883.4]
  wire  _T_15759; // @[Mux.scala 46:19:@12884.4]
  wire [7:0] _T_15760; // @[Mux.scala 46:16:@12885.4]
  wire  _T_15761; // @[Mux.scala 46:19:@12886.4]
  wire [7:0] _T_15762; // @[Mux.scala 46:16:@12887.4]
  wire  _T_15763; // @[Mux.scala 46:19:@12888.4]
  wire [7:0] _T_15764; // @[Mux.scala 46:16:@12889.4]
  wire  _T_15765; // @[Mux.scala 46:19:@12890.4]
  wire [7:0] _T_15766; // @[Mux.scala 46:16:@12891.4]
  wire  _T_15767; // @[Mux.scala 46:19:@12892.4]
  wire [7:0] _T_15768; // @[Mux.scala 46:16:@12893.4]
  wire  _T_15769; // @[Mux.scala 46:19:@12894.4]
  wire [7:0] _T_15770; // @[Mux.scala 46:16:@12895.4]
  wire  _T_15771; // @[Mux.scala 46:19:@12896.4]
  wire [7:0] _T_15772; // @[Mux.scala 46:16:@12897.4]
  wire  _T_15773; // @[Mux.scala 46:19:@12898.4]
  wire [7:0] _T_15774; // @[Mux.scala 46:16:@12899.4]
  wire  _T_15775; // @[Mux.scala 46:19:@12900.4]
  wire [7:0] _T_15776; // @[Mux.scala 46:16:@12901.4]
  wire  _T_15777; // @[Mux.scala 46:19:@12902.4]
  wire [7:0] _T_15778; // @[Mux.scala 46:16:@12903.4]
  wire  _T_15840; // @[Mux.scala 46:19:@12905.4]
  wire [7:0] _T_15841; // @[Mux.scala 46:16:@12906.4]
  wire  _T_15842; // @[Mux.scala 46:19:@12907.4]
  wire [7:0] _T_15843; // @[Mux.scala 46:16:@12908.4]
  wire  _T_15844; // @[Mux.scala 46:19:@12909.4]
  wire [7:0] _T_15845; // @[Mux.scala 46:16:@12910.4]
  wire  _T_15846; // @[Mux.scala 46:19:@12911.4]
  wire [7:0] _T_15847; // @[Mux.scala 46:16:@12912.4]
  wire  _T_15848; // @[Mux.scala 46:19:@12913.4]
  wire [7:0] _T_15849; // @[Mux.scala 46:16:@12914.4]
  wire  _T_15850; // @[Mux.scala 46:19:@12915.4]
  wire [7:0] _T_15851; // @[Mux.scala 46:16:@12916.4]
  wire  _T_15852; // @[Mux.scala 46:19:@12917.4]
  wire [7:0] _T_15853; // @[Mux.scala 46:16:@12918.4]
  wire  _T_15854; // @[Mux.scala 46:19:@12919.4]
  wire [7:0] _T_15855; // @[Mux.scala 46:16:@12920.4]
  wire  _T_15856; // @[Mux.scala 46:19:@12921.4]
  wire [7:0] _T_15857; // @[Mux.scala 46:16:@12922.4]
  wire  _T_15858; // @[Mux.scala 46:19:@12923.4]
  wire [7:0] _T_15859; // @[Mux.scala 46:16:@12924.4]
  wire  _T_15860; // @[Mux.scala 46:19:@12925.4]
  wire [7:0] _T_15861; // @[Mux.scala 46:16:@12926.4]
  wire  _T_15862; // @[Mux.scala 46:19:@12927.4]
  wire [7:0] _T_15863; // @[Mux.scala 46:16:@12928.4]
  wire  _T_15864; // @[Mux.scala 46:19:@12929.4]
  wire [7:0] _T_15865; // @[Mux.scala 46:16:@12930.4]
  wire  _T_15866; // @[Mux.scala 46:19:@12931.4]
  wire [7:0] _T_15867; // @[Mux.scala 46:16:@12932.4]
  wire  _T_15868; // @[Mux.scala 46:19:@12933.4]
  wire [7:0] _T_15869; // @[Mux.scala 46:16:@12934.4]
  wire  _T_15870; // @[Mux.scala 46:19:@12935.4]
  wire [7:0] _T_15871; // @[Mux.scala 46:16:@12936.4]
  wire  _T_15872; // @[Mux.scala 46:19:@12937.4]
  wire [7:0] _T_15873; // @[Mux.scala 46:16:@12938.4]
  wire  _T_15874; // @[Mux.scala 46:19:@12939.4]
  wire [7:0] _T_15875; // @[Mux.scala 46:16:@12940.4]
  wire  _T_15876; // @[Mux.scala 46:19:@12941.4]
  wire [7:0] _T_15877; // @[Mux.scala 46:16:@12942.4]
  wire  _T_15878; // @[Mux.scala 46:19:@12943.4]
  wire [7:0] _T_15879; // @[Mux.scala 46:16:@12944.4]
  wire  _T_15880; // @[Mux.scala 46:19:@12945.4]
  wire [7:0] _T_15881; // @[Mux.scala 46:16:@12946.4]
  wire  _T_15882; // @[Mux.scala 46:19:@12947.4]
  wire [7:0] _T_15883; // @[Mux.scala 46:16:@12948.4]
  wire  _T_15884; // @[Mux.scala 46:19:@12949.4]
  wire [7:0] _T_15885; // @[Mux.scala 46:16:@12950.4]
  wire  _T_15886; // @[Mux.scala 46:19:@12951.4]
  wire [7:0] _T_15887; // @[Mux.scala 46:16:@12952.4]
  wire  _T_15888; // @[Mux.scala 46:19:@12953.4]
  wire [7:0] _T_15889; // @[Mux.scala 46:16:@12954.4]
  wire  _T_15890; // @[Mux.scala 46:19:@12955.4]
  wire [7:0] _T_15891; // @[Mux.scala 46:16:@12956.4]
  wire  _T_15892; // @[Mux.scala 46:19:@12957.4]
  wire [7:0] _T_15893; // @[Mux.scala 46:16:@12958.4]
  wire  _T_15894; // @[Mux.scala 46:19:@12959.4]
  wire [7:0] _T_15895; // @[Mux.scala 46:16:@12960.4]
  wire  _T_15896; // @[Mux.scala 46:19:@12961.4]
  wire [7:0] _T_15897; // @[Mux.scala 46:16:@12962.4]
  wire  _T_15898; // @[Mux.scala 46:19:@12963.4]
  wire [7:0] _T_15899; // @[Mux.scala 46:16:@12964.4]
  wire  _T_15900; // @[Mux.scala 46:19:@12965.4]
  wire [7:0] _T_15901; // @[Mux.scala 46:16:@12966.4]
  wire  _T_15902; // @[Mux.scala 46:19:@12967.4]
  wire [7:0] _T_15903; // @[Mux.scala 46:16:@12968.4]
  wire  _T_15904; // @[Mux.scala 46:19:@12969.4]
  wire [7:0] _T_15905; // @[Mux.scala 46:16:@12970.4]
  wire  _T_15906; // @[Mux.scala 46:19:@12971.4]
  wire [7:0] _T_15907; // @[Mux.scala 46:16:@12972.4]
  wire  _T_15908; // @[Mux.scala 46:19:@12973.4]
  wire [7:0] _T_15909; // @[Mux.scala 46:16:@12974.4]
  wire  _T_15910; // @[Mux.scala 46:19:@12975.4]
  wire [7:0] _T_15911; // @[Mux.scala 46:16:@12976.4]
  wire  _T_15912; // @[Mux.scala 46:19:@12977.4]
  wire [7:0] _T_15913; // @[Mux.scala 46:16:@12978.4]
  wire  _T_15914; // @[Mux.scala 46:19:@12979.4]
  wire [7:0] _T_15915; // @[Mux.scala 46:16:@12980.4]
  wire  _T_15916; // @[Mux.scala 46:19:@12981.4]
  wire [7:0] _T_15917; // @[Mux.scala 46:16:@12982.4]
  wire  _T_15918; // @[Mux.scala 46:19:@12983.4]
  wire [7:0] _T_15919; // @[Mux.scala 46:16:@12984.4]
  wire  _T_15920; // @[Mux.scala 46:19:@12985.4]
  wire [7:0] _T_15921; // @[Mux.scala 46:16:@12986.4]
  wire  _T_15922; // @[Mux.scala 46:19:@12987.4]
  wire [7:0] _T_15923; // @[Mux.scala 46:16:@12988.4]
  wire  _T_15924; // @[Mux.scala 46:19:@12989.4]
  wire [7:0] _T_15925; // @[Mux.scala 46:16:@12990.4]
  wire  _T_15926; // @[Mux.scala 46:19:@12991.4]
  wire [7:0] _T_15927; // @[Mux.scala 46:16:@12992.4]
  wire  _T_15928; // @[Mux.scala 46:19:@12993.4]
  wire [7:0] _T_15929; // @[Mux.scala 46:16:@12994.4]
  wire  _T_15930; // @[Mux.scala 46:19:@12995.4]
  wire [7:0] _T_15931; // @[Mux.scala 46:16:@12996.4]
  wire  _T_15932; // @[Mux.scala 46:19:@12997.4]
  wire [7:0] _T_15933; // @[Mux.scala 46:16:@12998.4]
  wire  _T_15934; // @[Mux.scala 46:19:@12999.4]
  wire [7:0] _T_15935; // @[Mux.scala 46:16:@13000.4]
  wire  _T_15936; // @[Mux.scala 46:19:@13001.4]
  wire [7:0] _T_15937; // @[Mux.scala 46:16:@13002.4]
  wire  _T_15938; // @[Mux.scala 46:19:@13003.4]
  wire [7:0] _T_15939; // @[Mux.scala 46:16:@13004.4]
  wire  _T_15940; // @[Mux.scala 46:19:@13005.4]
  wire [7:0] _T_15941; // @[Mux.scala 46:16:@13006.4]
  wire  _T_15942; // @[Mux.scala 46:19:@13007.4]
  wire [7:0] _T_15943; // @[Mux.scala 46:16:@13008.4]
  wire  _T_15944; // @[Mux.scala 46:19:@13009.4]
  wire [7:0] _T_15945; // @[Mux.scala 46:16:@13010.4]
  wire  _T_15946; // @[Mux.scala 46:19:@13011.4]
  wire [7:0] _T_15947; // @[Mux.scala 46:16:@13012.4]
  wire  _T_15948; // @[Mux.scala 46:19:@13013.4]
  wire [7:0] _T_15949; // @[Mux.scala 46:16:@13014.4]
  wire  _T_15950; // @[Mux.scala 46:19:@13015.4]
  wire [7:0] _T_15951; // @[Mux.scala 46:16:@13016.4]
  wire  _T_15952; // @[Mux.scala 46:19:@13017.4]
  wire [7:0] _T_15953; // @[Mux.scala 46:16:@13018.4]
  wire  _T_15954; // @[Mux.scala 46:19:@13019.4]
  wire [7:0] _T_15955; // @[Mux.scala 46:16:@13020.4]
  wire  _T_15956; // @[Mux.scala 46:19:@13021.4]
  wire [7:0] _T_15957; // @[Mux.scala 46:16:@13022.4]
  wire  _T_15958; // @[Mux.scala 46:19:@13023.4]
  wire [7:0] _T_15959; // @[Mux.scala 46:16:@13024.4]
  wire  _T_16022; // @[Mux.scala 46:19:@13026.4]
  wire [7:0] _T_16023; // @[Mux.scala 46:16:@13027.4]
  wire  _T_16024; // @[Mux.scala 46:19:@13028.4]
  wire [7:0] _T_16025; // @[Mux.scala 46:16:@13029.4]
  wire  _T_16026; // @[Mux.scala 46:19:@13030.4]
  wire [7:0] _T_16027; // @[Mux.scala 46:16:@13031.4]
  wire  _T_16028; // @[Mux.scala 46:19:@13032.4]
  wire [7:0] _T_16029; // @[Mux.scala 46:16:@13033.4]
  wire  _T_16030; // @[Mux.scala 46:19:@13034.4]
  wire [7:0] _T_16031; // @[Mux.scala 46:16:@13035.4]
  wire  _T_16032; // @[Mux.scala 46:19:@13036.4]
  wire [7:0] _T_16033; // @[Mux.scala 46:16:@13037.4]
  wire  _T_16034; // @[Mux.scala 46:19:@13038.4]
  wire [7:0] _T_16035; // @[Mux.scala 46:16:@13039.4]
  wire  _T_16036; // @[Mux.scala 46:19:@13040.4]
  wire [7:0] _T_16037; // @[Mux.scala 46:16:@13041.4]
  wire  _T_16038; // @[Mux.scala 46:19:@13042.4]
  wire [7:0] _T_16039; // @[Mux.scala 46:16:@13043.4]
  wire  _T_16040; // @[Mux.scala 46:19:@13044.4]
  wire [7:0] _T_16041; // @[Mux.scala 46:16:@13045.4]
  wire  _T_16042; // @[Mux.scala 46:19:@13046.4]
  wire [7:0] _T_16043; // @[Mux.scala 46:16:@13047.4]
  wire  _T_16044; // @[Mux.scala 46:19:@13048.4]
  wire [7:0] _T_16045; // @[Mux.scala 46:16:@13049.4]
  wire  _T_16046; // @[Mux.scala 46:19:@13050.4]
  wire [7:0] _T_16047; // @[Mux.scala 46:16:@13051.4]
  wire  _T_16048; // @[Mux.scala 46:19:@13052.4]
  wire [7:0] _T_16049; // @[Mux.scala 46:16:@13053.4]
  wire  _T_16050; // @[Mux.scala 46:19:@13054.4]
  wire [7:0] _T_16051; // @[Mux.scala 46:16:@13055.4]
  wire  _T_16052; // @[Mux.scala 46:19:@13056.4]
  wire [7:0] _T_16053; // @[Mux.scala 46:16:@13057.4]
  wire  _T_16054; // @[Mux.scala 46:19:@13058.4]
  wire [7:0] _T_16055; // @[Mux.scala 46:16:@13059.4]
  wire  _T_16056; // @[Mux.scala 46:19:@13060.4]
  wire [7:0] _T_16057; // @[Mux.scala 46:16:@13061.4]
  wire  _T_16058; // @[Mux.scala 46:19:@13062.4]
  wire [7:0] _T_16059; // @[Mux.scala 46:16:@13063.4]
  wire  _T_16060; // @[Mux.scala 46:19:@13064.4]
  wire [7:0] _T_16061; // @[Mux.scala 46:16:@13065.4]
  wire  _T_16062; // @[Mux.scala 46:19:@13066.4]
  wire [7:0] _T_16063; // @[Mux.scala 46:16:@13067.4]
  wire  _T_16064; // @[Mux.scala 46:19:@13068.4]
  wire [7:0] _T_16065; // @[Mux.scala 46:16:@13069.4]
  wire  _T_16066; // @[Mux.scala 46:19:@13070.4]
  wire [7:0] _T_16067; // @[Mux.scala 46:16:@13071.4]
  wire  _T_16068; // @[Mux.scala 46:19:@13072.4]
  wire [7:0] _T_16069; // @[Mux.scala 46:16:@13073.4]
  wire  _T_16070; // @[Mux.scala 46:19:@13074.4]
  wire [7:0] _T_16071; // @[Mux.scala 46:16:@13075.4]
  wire  _T_16072; // @[Mux.scala 46:19:@13076.4]
  wire [7:0] _T_16073; // @[Mux.scala 46:16:@13077.4]
  wire  _T_16074; // @[Mux.scala 46:19:@13078.4]
  wire [7:0] _T_16075; // @[Mux.scala 46:16:@13079.4]
  wire  _T_16076; // @[Mux.scala 46:19:@13080.4]
  wire [7:0] _T_16077; // @[Mux.scala 46:16:@13081.4]
  wire  _T_16078; // @[Mux.scala 46:19:@13082.4]
  wire [7:0] _T_16079; // @[Mux.scala 46:16:@13083.4]
  wire  _T_16080; // @[Mux.scala 46:19:@13084.4]
  wire [7:0] _T_16081; // @[Mux.scala 46:16:@13085.4]
  wire  _T_16082; // @[Mux.scala 46:19:@13086.4]
  wire [7:0] _T_16083; // @[Mux.scala 46:16:@13087.4]
  wire  _T_16084; // @[Mux.scala 46:19:@13088.4]
  wire [7:0] _T_16085; // @[Mux.scala 46:16:@13089.4]
  wire  _T_16086; // @[Mux.scala 46:19:@13090.4]
  wire [7:0] _T_16087; // @[Mux.scala 46:16:@13091.4]
  wire  _T_16088; // @[Mux.scala 46:19:@13092.4]
  wire [7:0] _T_16089; // @[Mux.scala 46:16:@13093.4]
  wire  _T_16090; // @[Mux.scala 46:19:@13094.4]
  wire [7:0] _T_16091; // @[Mux.scala 46:16:@13095.4]
  wire  _T_16092; // @[Mux.scala 46:19:@13096.4]
  wire [7:0] _T_16093; // @[Mux.scala 46:16:@13097.4]
  wire  _T_16094; // @[Mux.scala 46:19:@13098.4]
  wire [7:0] _T_16095; // @[Mux.scala 46:16:@13099.4]
  wire  _T_16096; // @[Mux.scala 46:19:@13100.4]
  wire [7:0] _T_16097; // @[Mux.scala 46:16:@13101.4]
  wire  _T_16098; // @[Mux.scala 46:19:@13102.4]
  wire [7:0] _T_16099; // @[Mux.scala 46:16:@13103.4]
  wire  _T_16100; // @[Mux.scala 46:19:@13104.4]
  wire [7:0] _T_16101; // @[Mux.scala 46:16:@13105.4]
  wire  _T_16102; // @[Mux.scala 46:19:@13106.4]
  wire [7:0] _T_16103; // @[Mux.scala 46:16:@13107.4]
  wire  _T_16104; // @[Mux.scala 46:19:@13108.4]
  wire [7:0] _T_16105; // @[Mux.scala 46:16:@13109.4]
  wire  _T_16106; // @[Mux.scala 46:19:@13110.4]
  wire [7:0] _T_16107; // @[Mux.scala 46:16:@13111.4]
  wire  _T_16108; // @[Mux.scala 46:19:@13112.4]
  wire [7:0] _T_16109; // @[Mux.scala 46:16:@13113.4]
  wire  _T_16110; // @[Mux.scala 46:19:@13114.4]
  wire [7:0] _T_16111; // @[Mux.scala 46:16:@13115.4]
  wire  _T_16112; // @[Mux.scala 46:19:@13116.4]
  wire [7:0] _T_16113; // @[Mux.scala 46:16:@13117.4]
  wire  _T_16114; // @[Mux.scala 46:19:@13118.4]
  wire [7:0] _T_16115; // @[Mux.scala 46:16:@13119.4]
  wire  _T_16116; // @[Mux.scala 46:19:@13120.4]
  wire [7:0] _T_16117; // @[Mux.scala 46:16:@13121.4]
  wire  _T_16118; // @[Mux.scala 46:19:@13122.4]
  wire [7:0] _T_16119; // @[Mux.scala 46:16:@13123.4]
  wire  _T_16120; // @[Mux.scala 46:19:@13124.4]
  wire [7:0] _T_16121; // @[Mux.scala 46:16:@13125.4]
  wire  _T_16122; // @[Mux.scala 46:19:@13126.4]
  wire [7:0] _T_16123; // @[Mux.scala 46:16:@13127.4]
  wire  _T_16124; // @[Mux.scala 46:19:@13128.4]
  wire [7:0] _T_16125; // @[Mux.scala 46:16:@13129.4]
  wire  _T_16126; // @[Mux.scala 46:19:@13130.4]
  wire [7:0] _T_16127; // @[Mux.scala 46:16:@13131.4]
  wire  _T_16128; // @[Mux.scala 46:19:@13132.4]
  wire [7:0] _T_16129; // @[Mux.scala 46:16:@13133.4]
  wire  _T_16130; // @[Mux.scala 46:19:@13134.4]
  wire [7:0] _T_16131; // @[Mux.scala 46:16:@13135.4]
  wire  _T_16132; // @[Mux.scala 46:19:@13136.4]
  wire [7:0] _T_16133; // @[Mux.scala 46:16:@13137.4]
  wire  _T_16134; // @[Mux.scala 46:19:@13138.4]
  wire [7:0] _T_16135; // @[Mux.scala 46:16:@13139.4]
  wire  _T_16136; // @[Mux.scala 46:19:@13140.4]
  wire [7:0] _T_16137; // @[Mux.scala 46:16:@13141.4]
  wire  _T_16138; // @[Mux.scala 46:19:@13142.4]
  wire [7:0] _T_16139; // @[Mux.scala 46:16:@13143.4]
  wire  _T_16140; // @[Mux.scala 46:19:@13144.4]
  wire [7:0] _T_16141; // @[Mux.scala 46:16:@13145.4]
  wire  _T_16142; // @[Mux.scala 46:19:@13146.4]
  wire [7:0] _T_16143; // @[Mux.scala 46:16:@13147.4]
  wire  _T_16207; // @[Mux.scala 46:19:@13149.4]
  wire [7:0] _T_16208; // @[Mux.scala 46:16:@13150.4]
  wire  _T_16209; // @[Mux.scala 46:19:@13151.4]
  wire [7:0] _T_16210; // @[Mux.scala 46:16:@13152.4]
  wire  _T_16211; // @[Mux.scala 46:19:@13153.4]
  wire [7:0] _T_16212; // @[Mux.scala 46:16:@13154.4]
  wire  _T_16213; // @[Mux.scala 46:19:@13155.4]
  wire [7:0] _T_16214; // @[Mux.scala 46:16:@13156.4]
  wire  _T_16215; // @[Mux.scala 46:19:@13157.4]
  wire [7:0] _T_16216; // @[Mux.scala 46:16:@13158.4]
  wire  _T_16217; // @[Mux.scala 46:19:@13159.4]
  wire [7:0] _T_16218; // @[Mux.scala 46:16:@13160.4]
  wire  _T_16219; // @[Mux.scala 46:19:@13161.4]
  wire [7:0] _T_16220; // @[Mux.scala 46:16:@13162.4]
  wire  _T_16221; // @[Mux.scala 46:19:@13163.4]
  wire [7:0] _T_16222; // @[Mux.scala 46:16:@13164.4]
  wire  _T_16223; // @[Mux.scala 46:19:@13165.4]
  wire [7:0] _T_16224; // @[Mux.scala 46:16:@13166.4]
  wire  _T_16225; // @[Mux.scala 46:19:@13167.4]
  wire [7:0] _T_16226; // @[Mux.scala 46:16:@13168.4]
  wire  _T_16227; // @[Mux.scala 46:19:@13169.4]
  wire [7:0] _T_16228; // @[Mux.scala 46:16:@13170.4]
  wire  _T_16229; // @[Mux.scala 46:19:@13171.4]
  wire [7:0] _T_16230; // @[Mux.scala 46:16:@13172.4]
  wire  _T_16231; // @[Mux.scala 46:19:@13173.4]
  wire [7:0] _T_16232; // @[Mux.scala 46:16:@13174.4]
  wire  _T_16233; // @[Mux.scala 46:19:@13175.4]
  wire [7:0] _T_16234; // @[Mux.scala 46:16:@13176.4]
  wire  _T_16235; // @[Mux.scala 46:19:@13177.4]
  wire [7:0] _T_16236; // @[Mux.scala 46:16:@13178.4]
  wire  _T_16237; // @[Mux.scala 46:19:@13179.4]
  wire [7:0] _T_16238; // @[Mux.scala 46:16:@13180.4]
  wire  _T_16239; // @[Mux.scala 46:19:@13181.4]
  wire [7:0] _T_16240; // @[Mux.scala 46:16:@13182.4]
  wire  _T_16241; // @[Mux.scala 46:19:@13183.4]
  wire [7:0] _T_16242; // @[Mux.scala 46:16:@13184.4]
  wire  _T_16243; // @[Mux.scala 46:19:@13185.4]
  wire [7:0] _T_16244; // @[Mux.scala 46:16:@13186.4]
  wire  _T_16245; // @[Mux.scala 46:19:@13187.4]
  wire [7:0] _T_16246; // @[Mux.scala 46:16:@13188.4]
  wire  _T_16247; // @[Mux.scala 46:19:@13189.4]
  wire [7:0] _T_16248; // @[Mux.scala 46:16:@13190.4]
  wire  _T_16249; // @[Mux.scala 46:19:@13191.4]
  wire [7:0] _T_16250; // @[Mux.scala 46:16:@13192.4]
  wire  _T_16251; // @[Mux.scala 46:19:@13193.4]
  wire [7:0] _T_16252; // @[Mux.scala 46:16:@13194.4]
  wire  _T_16253; // @[Mux.scala 46:19:@13195.4]
  wire [7:0] _T_16254; // @[Mux.scala 46:16:@13196.4]
  wire  _T_16255; // @[Mux.scala 46:19:@13197.4]
  wire [7:0] _T_16256; // @[Mux.scala 46:16:@13198.4]
  wire  _T_16257; // @[Mux.scala 46:19:@13199.4]
  wire [7:0] _T_16258; // @[Mux.scala 46:16:@13200.4]
  wire  _T_16259; // @[Mux.scala 46:19:@13201.4]
  wire [7:0] _T_16260; // @[Mux.scala 46:16:@13202.4]
  wire  _T_16261; // @[Mux.scala 46:19:@13203.4]
  wire [7:0] _T_16262; // @[Mux.scala 46:16:@13204.4]
  wire  _T_16263; // @[Mux.scala 46:19:@13205.4]
  wire [7:0] _T_16264; // @[Mux.scala 46:16:@13206.4]
  wire  _T_16265; // @[Mux.scala 46:19:@13207.4]
  wire [7:0] _T_16266; // @[Mux.scala 46:16:@13208.4]
  wire  _T_16267; // @[Mux.scala 46:19:@13209.4]
  wire [7:0] _T_16268; // @[Mux.scala 46:16:@13210.4]
  wire  _T_16269; // @[Mux.scala 46:19:@13211.4]
  wire [7:0] _T_16270; // @[Mux.scala 46:16:@13212.4]
  wire  _T_16271; // @[Mux.scala 46:19:@13213.4]
  wire [7:0] _T_16272; // @[Mux.scala 46:16:@13214.4]
  wire  _T_16273; // @[Mux.scala 46:19:@13215.4]
  wire [7:0] _T_16274; // @[Mux.scala 46:16:@13216.4]
  wire  _T_16275; // @[Mux.scala 46:19:@13217.4]
  wire [7:0] _T_16276; // @[Mux.scala 46:16:@13218.4]
  wire  _T_16277; // @[Mux.scala 46:19:@13219.4]
  wire [7:0] _T_16278; // @[Mux.scala 46:16:@13220.4]
  wire  _T_16279; // @[Mux.scala 46:19:@13221.4]
  wire [7:0] _T_16280; // @[Mux.scala 46:16:@13222.4]
  wire  _T_16281; // @[Mux.scala 46:19:@13223.4]
  wire [7:0] _T_16282; // @[Mux.scala 46:16:@13224.4]
  wire  _T_16283; // @[Mux.scala 46:19:@13225.4]
  wire [7:0] _T_16284; // @[Mux.scala 46:16:@13226.4]
  wire  _T_16285; // @[Mux.scala 46:19:@13227.4]
  wire [7:0] _T_16286; // @[Mux.scala 46:16:@13228.4]
  wire  _T_16287; // @[Mux.scala 46:19:@13229.4]
  wire [7:0] _T_16288; // @[Mux.scala 46:16:@13230.4]
  wire  _T_16289; // @[Mux.scala 46:19:@13231.4]
  wire [7:0] _T_16290; // @[Mux.scala 46:16:@13232.4]
  wire  _T_16291; // @[Mux.scala 46:19:@13233.4]
  wire [7:0] _T_16292; // @[Mux.scala 46:16:@13234.4]
  wire  _T_16293; // @[Mux.scala 46:19:@13235.4]
  wire [7:0] _T_16294; // @[Mux.scala 46:16:@13236.4]
  wire  _T_16295; // @[Mux.scala 46:19:@13237.4]
  wire [7:0] _T_16296; // @[Mux.scala 46:16:@13238.4]
  wire  _T_16297; // @[Mux.scala 46:19:@13239.4]
  wire [7:0] _T_16298; // @[Mux.scala 46:16:@13240.4]
  wire  _T_16299; // @[Mux.scala 46:19:@13241.4]
  wire [7:0] _T_16300; // @[Mux.scala 46:16:@13242.4]
  wire  _T_16301; // @[Mux.scala 46:19:@13243.4]
  wire [7:0] _T_16302; // @[Mux.scala 46:16:@13244.4]
  wire  _T_16303; // @[Mux.scala 46:19:@13245.4]
  wire [7:0] _T_16304; // @[Mux.scala 46:16:@13246.4]
  wire  _T_16305; // @[Mux.scala 46:19:@13247.4]
  wire [7:0] _T_16306; // @[Mux.scala 46:16:@13248.4]
  wire  _T_16307; // @[Mux.scala 46:19:@13249.4]
  wire [7:0] _T_16308; // @[Mux.scala 46:16:@13250.4]
  wire  _T_16309; // @[Mux.scala 46:19:@13251.4]
  wire [7:0] _T_16310; // @[Mux.scala 46:16:@13252.4]
  wire  _T_16311; // @[Mux.scala 46:19:@13253.4]
  wire [7:0] _T_16312; // @[Mux.scala 46:16:@13254.4]
  wire  _T_16313; // @[Mux.scala 46:19:@13255.4]
  wire [7:0] _T_16314; // @[Mux.scala 46:16:@13256.4]
  wire  _T_16315; // @[Mux.scala 46:19:@13257.4]
  wire [7:0] _T_16316; // @[Mux.scala 46:16:@13258.4]
  wire  _T_16317; // @[Mux.scala 46:19:@13259.4]
  wire [7:0] _T_16318; // @[Mux.scala 46:16:@13260.4]
  wire  _T_16319; // @[Mux.scala 46:19:@13261.4]
  wire [7:0] _T_16320; // @[Mux.scala 46:16:@13262.4]
  wire  _T_16321; // @[Mux.scala 46:19:@13263.4]
  wire [7:0] _T_16322; // @[Mux.scala 46:16:@13264.4]
  wire  _T_16323; // @[Mux.scala 46:19:@13265.4]
  wire [7:0] _T_16324; // @[Mux.scala 46:16:@13266.4]
  wire  _T_16325; // @[Mux.scala 46:19:@13267.4]
  wire [7:0] _T_16326; // @[Mux.scala 46:16:@13268.4]
  wire  _T_16327; // @[Mux.scala 46:19:@13269.4]
  wire [7:0] _T_16328; // @[Mux.scala 46:16:@13270.4]
  wire  _T_16329; // @[Mux.scala 46:19:@13271.4]
  wire [7:0] _T_16330; // @[Mux.scala 46:16:@13272.4]
  wire  _T_16395; // @[Mux.scala 46:19:@13274.4]
  wire [7:0] _T_16396; // @[Mux.scala 46:16:@13275.4]
  wire  _T_16397; // @[Mux.scala 46:19:@13276.4]
  wire [7:0] _T_16398; // @[Mux.scala 46:16:@13277.4]
  wire  _T_16399; // @[Mux.scala 46:19:@13278.4]
  wire [7:0] _T_16400; // @[Mux.scala 46:16:@13279.4]
  wire  _T_16401; // @[Mux.scala 46:19:@13280.4]
  wire [7:0] _T_16402; // @[Mux.scala 46:16:@13281.4]
  wire  _T_16403; // @[Mux.scala 46:19:@13282.4]
  wire [7:0] _T_16404; // @[Mux.scala 46:16:@13283.4]
  wire  _T_16405; // @[Mux.scala 46:19:@13284.4]
  wire [7:0] _T_16406; // @[Mux.scala 46:16:@13285.4]
  wire  _T_16407; // @[Mux.scala 46:19:@13286.4]
  wire [7:0] _T_16408; // @[Mux.scala 46:16:@13287.4]
  wire  _T_16409; // @[Mux.scala 46:19:@13288.4]
  wire [7:0] _T_16410; // @[Mux.scala 46:16:@13289.4]
  wire  _T_16411; // @[Mux.scala 46:19:@13290.4]
  wire [7:0] _T_16412; // @[Mux.scala 46:16:@13291.4]
  wire  _T_16413; // @[Mux.scala 46:19:@13292.4]
  wire [7:0] _T_16414; // @[Mux.scala 46:16:@13293.4]
  wire  _T_16415; // @[Mux.scala 46:19:@13294.4]
  wire [7:0] _T_16416; // @[Mux.scala 46:16:@13295.4]
  wire  _T_16417; // @[Mux.scala 46:19:@13296.4]
  wire [7:0] _T_16418; // @[Mux.scala 46:16:@13297.4]
  wire  _T_16419; // @[Mux.scala 46:19:@13298.4]
  wire [7:0] _T_16420; // @[Mux.scala 46:16:@13299.4]
  wire  _T_16421; // @[Mux.scala 46:19:@13300.4]
  wire [7:0] _T_16422; // @[Mux.scala 46:16:@13301.4]
  wire  _T_16423; // @[Mux.scala 46:19:@13302.4]
  wire [7:0] _T_16424; // @[Mux.scala 46:16:@13303.4]
  wire  _T_16425; // @[Mux.scala 46:19:@13304.4]
  wire [7:0] _T_16426; // @[Mux.scala 46:16:@13305.4]
  wire  _T_16427; // @[Mux.scala 46:19:@13306.4]
  wire [7:0] _T_16428; // @[Mux.scala 46:16:@13307.4]
  wire  _T_16429; // @[Mux.scala 46:19:@13308.4]
  wire [7:0] _T_16430; // @[Mux.scala 46:16:@13309.4]
  wire  _T_16431; // @[Mux.scala 46:19:@13310.4]
  wire [7:0] _T_16432; // @[Mux.scala 46:16:@13311.4]
  wire  _T_16433; // @[Mux.scala 46:19:@13312.4]
  wire [7:0] _T_16434; // @[Mux.scala 46:16:@13313.4]
  wire  _T_16435; // @[Mux.scala 46:19:@13314.4]
  wire [7:0] _T_16436; // @[Mux.scala 46:16:@13315.4]
  wire  _T_16437; // @[Mux.scala 46:19:@13316.4]
  wire [7:0] _T_16438; // @[Mux.scala 46:16:@13317.4]
  wire  _T_16439; // @[Mux.scala 46:19:@13318.4]
  wire [7:0] _T_16440; // @[Mux.scala 46:16:@13319.4]
  wire  _T_16441; // @[Mux.scala 46:19:@13320.4]
  wire [7:0] _T_16442; // @[Mux.scala 46:16:@13321.4]
  wire  _T_16443; // @[Mux.scala 46:19:@13322.4]
  wire [7:0] _T_16444; // @[Mux.scala 46:16:@13323.4]
  wire  _T_16445; // @[Mux.scala 46:19:@13324.4]
  wire [7:0] _T_16446; // @[Mux.scala 46:16:@13325.4]
  wire  _T_16447; // @[Mux.scala 46:19:@13326.4]
  wire [7:0] _T_16448; // @[Mux.scala 46:16:@13327.4]
  wire  _T_16449; // @[Mux.scala 46:19:@13328.4]
  wire [7:0] _T_16450; // @[Mux.scala 46:16:@13329.4]
  wire  _T_16451; // @[Mux.scala 46:19:@13330.4]
  wire [7:0] _T_16452; // @[Mux.scala 46:16:@13331.4]
  wire  _T_16453; // @[Mux.scala 46:19:@13332.4]
  wire [7:0] _T_16454; // @[Mux.scala 46:16:@13333.4]
  wire  _T_16455; // @[Mux.scala 46:19:@13334.4]
  wire [7:0] _T_16456; // @[Mux.scala 46:16:@13335.4]
  wire  _T_16457; // @[Mux.scala 46:19:@13336.4]
  wire [7:0] _T_16458; // @[Mux.scala 46:16:@13337.4]
  wire  _T_16459; // @[Mux.scala 46:19:@13338.4]
  wire [7:0] _T_16460; // @[Mux.scala 46:16:@13339.4]
  wire  _T_16461; // @[Mux.scala 46:19:@13340.4]
  wire [7:0] _T_16462; // @[Mux.scala 46:16:@13341.4]
  wire  _T_16463; // @[Mux.scala 46:19:@13342.4]
  wire [7:0] _T_16464; // @[Mux.scala 46:16:@13343.4]
  wire  _T_16465; // @[Mux.scala 46:19:@13344.4]
  wire [7:0] _T_16466; // @[Mux.scala 46:16:@13345.4]
  wire  _T_16467; // @[Mux.scala 46:19:@13346.4]
  wire [7:0] _T_16468; // @[Mux.scala 46:16:@13347.4]
  wire  _T_16469; // @[Mux.scala 46:19:@13348.4]
  wire [7:0] _T_16470; // @[Mux.scala 46:16:@13349.4]
  wire  _T_16471; // @[Mux.scala 46:19:@13350.4]
  wire [7:0] _T_16472; // @[Mux.scala 46:16:@13351.4]
  wire  _T_16473; // @[Mux.scala 46:19:@13352.4]
  wire [7:0] _T_16474; // @[Mux.scala 46:16:@13353.4]
  wire  _T_16475; // @[Mux.scala 46:19:@13354.4]
  wire [7:0] _T_16476; // @[Mux.scala 46:16:@13355.4]
  wire  _T_16477; // @[Mux.scala 46:19:@13356.4]
  wire [7:0] _T_16478; // @[Mux.scala 46:16:@13357.4]
  wire  _T_16479; // @[Mux.scala 46:19:@13358.4]
  wire [7:0] _T_16480; // @[Mux.scala 46:16:@13359.4]
  wire  _T_16481; // @[Mux.scala 46:19:@13360.4]
  wire [7:0] _T_16482; // @[Mux.scala 46:16:@13361.4]
  wire  _T_16483; // @[Mux.scala 46:19:@13362.4]
  wire [7:0] _T_16484; // @[Mux.scala 46:16:@13363.4]
  wire  _T_16485; // @[Mux.scala 46:19:@13364.4]
  wire [7:0] _T_16486; // @[Mux.scala 46:16:@13365.4]
  wire  _T_16487; // @[Mux.scala 46:19:@13366.4]
  wire [7:0] _T_16488; // @[Mux.scala 46:16:@13367.4]
  wire  _T_16489; // @[Mux.scala 46:19:@13368.4]
  wire [7:0] _T_16490; // @[Mux.scala 46:16:@13369.4]
  wire  _T_16491; // @[Mux.scala 46:19:@13370.4]
  wire [7:0] _T_16492; // @[Mux.scala 46:16:@13371.4]
  wire  _T_16493; // @[Mux.scala 46:19:@13372.4]
  wire [7:0] _T_16494; // @[Mux.scala 46:16:@13373.4]
  wire  _T_16495; // @[Mux.scala 46:19:@13374.4]
  wire [7:0] _T_16496; // @[Mux.scala 46:16:@13375.4]
  wire  _T_16497; // @[Mux.scala 46:19:@13376.4]
  wire [7:0] _T_16498; // @[Mux.scala 46:16:@13377.4]
  wire  _T_16499; // @[Mux.scala 46:19:@13378.4]
  wire [7:0] _T_16500; // @[Mux.scala 46:16:@13379.4]
  wire  _T_16501; // @[Mux.scala 46:19:@13380.4]
  wire [7:0] _T_16502; // @[Mux.scala 46:16:@13381.4]
  wire  _T_16503; // @[Mux.scala 46:19:@13382.4]
  wire [7:0] _T_16504; // @[Mux.scala 46:16:@13383.4]
  wire  _T_16505; // @[Mux.scala 46:19:@13384.4]
  wire [7:0] _T_16506; // @[Mux.scala 46:16:@13385.4]
  wire  _T_16507; // @[Mux.scala 46:19:@13386.4]
  wire [7:0] _T_16508; // @[Mux.scala 46:16:@13387.4]
  wire  _T_16509; // @[Mux.scala 46:19:@13388.4]
  wire [7:0] _T_16510; // @[Mux.scala 46:16:@13389.4]
  wire  _T_16511; // @[Mux.scala 46:19:@13390.4]
  wire [7:0] _T_16512; // @[Mux.scala 46:16:@13391.4]
  wire  _T_16513; // @[Mux.scala 46:19:@13392.4]
  wire [7:0] _T_16514; // @[Mux.scala 46:16:@13393.4]
  wire  _T_16515; // @[Mux.scala 46:19:@13394.4]
  wire [7:0] _T_16516; // @[Mux.scala 46:16:@13395.4]
  wire  _T_16517; // @[Mux.scala 46:19:@13396.4]
  wire [7:0] _T_16518; // @[Mux.scala 46:16:@13397.4]
  wire  _T_16519; // @[Mux.scala 46:19:@13398.4]
  wire [7:0] _T_16520; // @[Mux.scala 46:16:@13399.4]
  wire  _T_16586; // @[Mux.scala 46:19:@13401.4]
  wire [7:0] _T_16587; // @[Mux.scala 46:16:@13402.4]
  wire  _T_16588; // @[Mux.scala 46:19:@13403.4]
  wire [7:0] _T_16589; // @[Mux.scala 46:16:@13404.4]
  wire  _T_16590; // @[Mux.scala 46:19:@13405.4]
  wire [7:0] _T_16591; // @[Mux.scala 46:16:@13406.4]
  wire  _T_16592; // @[Mux.scala 46:19:@13407.4]
  wire [7:0] _T_16593; // @[Mux.scala 46:16:@13408.4]
  wire  _T_16594; // @[Mux.scala 46:19:@13409.4]
  wire [7:0] _T_16595; // @[Mux.scala 46:16:@13410.4]
  wire  _T_16596; // @[Mux.scala 46:19:@13411.4]
  wire [7:0] _T_16597; // @[Mux.scala 46:16:@13412.4]
  wire  _T_16598; // @[Mux.scala 46:19:@13413.4]
  wire [7:0] _T_16599; // @[Mux.scala 46:16:@13414.4]
  wire  _T_16600; // @[Mux.scala 46:19:@13415.4]
  wire [7:0] _T_16601; // @[Mux.scala 46:16:@13416.4]
  wire  _T_16602; // @[Mux.scala 46:19:@13417.4]
  wire [7:0] _T_16603; // @[Mux.scala 46:16:@13418.4]
  wire  _T_16604; // @[Mux.scala 46:19:@13419.4]
  wire [7:0] _T_16605; // @[Mux.scala 46:16:@13420.4]
  wire  _T_16606; // @[Mux.scala 46:19:@13421.4]
  wire [7:0] _T_16607; // @[Mux.scala 46:16:@13422.4]
  wire  _T_16608; // @[Mux.scala 46:19:@13423.4]
  wire [7:0] _T_16609; // @[Mux.scala 46:16:@13424.4]
  wire  _T_16610; // @[Mux.scala 46:19:@13425.4]
  wire [7:0] _T_16611; // @[Mux.scala 46:16:@13426.4]
  wire  _T_16612; // @[Mux.scala 46:19:@13427.4]
  wire [7:0] _T_16613; // @[Mux.scala 46:16:@13428.4]
  wire  _T_16614; // @[Mux.scala 46:19:@13429.4]
  wire [7:0] _T_16615; // @[Mux.scala 46:16:@13430.4]
  wire  _T_16616; // @[Mux.scala 46:19:@13431.4]
  wire [7:0] _T_16617; // @[Mux.scala 46:16:@13432.4]
  wire  _T_16618; // @[Mux.scala 46:19:@13433.4]
  wire [7:0] _T_16619; // @[Mux.scala 46:16:@13434.4]
  wire  _T_16620; // @[Mux.scala 46:19:@13435.4]
  wire [7:0] _T_16621; // @[Mux.scala 46:16:@13436.4]
  wire  _T_16622; // @[Mux.scala 46:19:@13437.4]
  wire [7:0] _T_16623; // @[Mux.scala 46:16:@13438.4]
  wire  _T_16624; // @[Mux.scala 46:19:@13439.4]
  wire [7:0] _T_16625; // @[Mux.scala 46:16:@13440.4]
  wire  _T_16626; // @[Mux.scala 46:19:@13441.4]
  wire [7:0] _T_16627; // @[Mux.scala 46:16:@13442.4]
  wire  _T_16628; // @[Mux.scala 46:19:@13443.4]
  wire [7:0] _T_16629; // @[Mux.scala 46:16:@13444.4]
  wire  _T_16630; // @[Mux.scala 46:19:@13445.4]
  wire [7:0] _T_16631; // @[Mux.scala 46:16:@13446.4]
  wire  _T_16632; // @[Mux.scala 46:19:@13447.4]
  wire [7:0] _T_16633; // @[Mux.scala 46:16:@13448.4]
  wire  _T_16634; // @[Mux.scala 46:19:@13449.4]
  wire [7:0] _T_16635; // @[Mux.scala 46:16:@13450.4]
  wire  _T_16636; // @[Mux.scala 46:19:@13451.4]
  wire [7:0] _T_16637; // @[Mux.scala 46:16:@13452.4]
  wire  _T_16638; // @[Mux.scala 46:19:@13453.4]
  wire [7:0] _T_16639; // @[Mux.scala 46:16:@13454.4]
  wire  _T_16640; // @[Mux.scala 46:19:@13455.4]
  wire [7:0] _T_16641; // @[Mux.scala 46:16:@13456.4]
  wire  _T_16642; // @[Mux.scala 46:19:@13457.4]
  wire [7:0] _T_16643; // @[Mux.scala 46:16:@13458.4]
  wire  _T_16644; // @[Mux.scala 46:19:@13459.4]
  wire [7:0] _T_16645; // @[Mux.scala 46:16:@13460.4]
  wire  _T_16646; // @[Mux.scala 46:19:@13461.4]
  wire [7:0] _T_16647; // @[Mux.scala 46:16:@13462.4]
  wire  _T_16648; // @[Mux.scala 46:19:@13463.4]
  wire [7:0] _T_16649; // @[Mux.scala 46:16:@13464.4]
  wire  _T_16650; // @[Mux.scala 46:19:@13465.4]
  wire [7:0] _T_16651; // @[Mux.scala 46:16:@13466.4]
  wire  _T_16652; // @[Mux.scala 46:19:@13467.4]
  wire [7:0] _T_16653; // @[Mux.scala 46:16:@13468.4]
  wire  _T_16654; // @[Mux.scala 46:19:@13469.4]
  wire [7:0] _T_16655; // @[Mux.scala 46:16:@13470.4]
  wire  _T_16656; // @[Mux.scala 46:19:@13471.4]
  wire [7:0] _T_16657; // @[Mux.scala 46:16:@13472.4]
  wire  _T_16658; // @[Mux.scala 46:19:@13473.4]
  wire [7:0] _T_16659; // @[Mux.scala 46:16:@13474.4]
  wire  _T_16660; // @[Mux.scala 46:19:@13475.4]
  wire [7:0] _T_16661; // @[Mux.scala 46:16:@13476.4]
  wire  _T_16662; // @[Mux.scala 46:19:@13477.4]
  wire [7:0] _T_16663; // @[Mux.scala 46:16:@13478.4]
  wire  _T_16664; // @[Mux.scala 46:19:@13479.4]
  wire [7:0] _T_16665; // @[Mux.scala 46:16:@13480.4]
  wire  _T_16666; // @[Mux.scala 46:19:@13481.4]
  wire [7:0] _T_16667; // @[Mux.scala 46:16:@13482.4]
  wire  _T_16668; // @[Mux.scala 46:19:@13483.4]
  wire [7:0] _T_16669; // @[Mux.scala 46:16:@13484.4]
  wire  _T_16670; // @[Mux.scala 46:19:@13485.4]
  wire [7:0] _T_16671; // @[Mux.scala 46:16:@13486.4]
  wire  _T_16672; // @[Mux.scala 46:19:@13487.4]
  wire [7:0] _T_16673; // @[Mux.scala 46:16:@13488.4]
  wire  _T_16674; // @[Mux.scala 46:19:@13489.4]
  wire [7:0] _T_16675; // @[Mux.scala 46:16:@13490.4]
  wire  _T_16676; // @[Mux.scala 46:19:@13491.4]
  wire [7:0] _T_16677; // @[Mux.scala 46:16:@13492.4]
  wire  _T_16678; // @[Mux.scala 46:19:@13493.4]
  wire [7:0] _T_16679; // @[Mux.scala 46:16:@13494.4]
  wire  _T_16680; // @[Mux.scala 46:19:@13495.4]
  wire [7:0] _T_16681; // @[Mux.scala 46:16:@13496.4]
  wire  _T_16682; // @[Mux.scala 46:19:@13497.4]
  wire [7:0] _T_16683; // @[Mux.scala 46:16:@13498.4]
  wire  _T_16684; // @[Mux.scala 46:19:@13499.4]
  wire [7:0] _T_16685; // @[Mux.scala 46:16:@13500.4]
  wire  _T_16686; // @[Mux.scala 46:19:@13501.4]
  wire [7:0] _T_16687; // @[Mux.scala 46:16:@13502.4]
  wire  _T_16688; // @[Mux.scala 46:19:@13503.4]
  wire [7:0] _T_16689; // @[Mux.scala 46:16:@13504.4]
  wire  _T_16690; // @[Mux.scala 46:19:@13505.4]
  wire [7:0] _T_16691; // @[Mux.scala 46:16:@13506.4]
  wire  _T_16692; // @[Mux.scala 46:19:@13507.4]
  wire [7:0] _T_16693; // @[Mux.scala 46:16:@13508.4]
  wire  _T_16694; // @[Mux.scala 46:19:@13509.4]
  wire [7:0] _T_16695; // @[Mux.scala 46:16:@13510.4]
  wire  _T_16696; // @[Mux.scala 46:19:@13511.4]
  wire [7:0] _T_16697; // @[Mux.scala 46:16:@13512.4]
  wire  _T_16698; // @[Mux.scala 46:19:@13513.4]
  wire [7:0] _T_16699; // @[Mux.scala 46:16:@13514.4]
  wire  _T_16700; // @[Mux.scala 46:19:@13515.4]
  wire [7:0] _T_16701; // @[Mux.scala 46:16:@13516.4]
  wire  _T_16702; // @[Mux.scala 46:19:@13517.4]
  wire [7:0] _T_16703; // @[Mux.scala 46:16:@13518.4]
  wire  _T_16704; // @[Mux.scala 46:19:@13519.4]
  wire [7:0] _T_16705; // @[Mux.scala 46:16:@13520.4]
  wire  _T_16706; // @[Mux.scala 46:19:@13521.4]
  wire [7:0] _T_16707; // @[Mux.scala 46:16:@13522.4]
  wire  _T_16708; // @[Mux.scala 46:19:@13523.4]
  wire [7:0] _T_16709; // @[Mux.scala 46:16:@13524.4]
  wire  _T_16710; // @[Mux.scala 46:19:@13525.4]
  wire [7:0] _T_16711; // @[Mux.scala 46:16:@13526.4]
  wire  _T_16712; // @[Mux.scala 46:19:@13527.4]
  wire [7:0] _T_16713; // @[Mux.scala 46:16:@13528.4]
  reg  _T_16716; // @[NV_NVDLA_CSC_WL_dec.scala 119:27:@13530.4]
  reg [31:0] _RAND_225;
  reg  _T_16855_0; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_226;
  reg  _T_16855_1; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_227;
  reg  _T_16855_2; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_228;
  reg  _T_16855_3; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_229;
  reg  _T_16855_4; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_230;
  reg  _T_16855_5; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_231;
  reg  _T_16855_6; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_232;
  reg  _T_16855_7; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_233;
  reg  _T_16855_8; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_234;
  reg  _T_16855_9; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_235;
  reg  _T_16855_10; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_236;
  reg  _T_16855_11; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_237;
  reg  _T_16855_12; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_238;
  reg  _T_16855_13; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_239;
  reg  _T_16855_14; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_240;
  reg  _T_16855_15; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_241;
  reg  _T_16855_16; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_242;
  reg  _T_16855_17; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_243;
  reg  _T_16855_18; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_244;
  reg  _T_16855_19; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_245;
  reg  _T_16855_20; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_246;
  reg  _T_16855_21; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_247;
  reg  _T_16855_22; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_248;
  reg  _T_16855_23; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_249;
  reg  _T_16855_24; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_250;
  reg  _T_16855_25; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_251;
  reg  _T_16855_26; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_252;
  reg  _T_16855_27; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_253;
  reg  _T_16855_28; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_254;
  reg  _T_16855_29; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_255;
  reg  _T_16855_30; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_256;
  reg  _T_16855_31; // @[NV_NVDLA_CSC_WL_dec.scala 120:25:@13564.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_16959_0; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_16959_1; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_16959_2; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_16959_3; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_16959_4; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_16959_5; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_16959_6; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_16959_7; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_16959_8; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_16959_9; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_16959_10; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_16959_11; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_16959_12; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_16959_13; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_16959_14; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_16959_15; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_16959_16; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_16959_17; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_16959_18; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_16959_19; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_16959_20; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_16959_21; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_16959_22; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_16959_23; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_281;
  reg [7:0] _T_16959_24; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_282;
  reg [7:0] _T_16959_25; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_283;
  reg [7:0] _T_16959_26; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_284;
  reg [7:0] _T_16959_27; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_285;
  reg [7:0] _T_16959_28; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_286;
  reg [7:0] _T_16959_29; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_287;
  reg [7:0] _T_16959_30; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_288;
  reg [7:0] _T_16959_31; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_289;
  reg [7:0] _T_16959_32; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_290;
  reg [7:0] _T_16959_33; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_291;
  reg [7:0] _T_16959_34; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_292;
  reg [7:0] _T_16959_35; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_293;
  reg [7:0] _T_16959_36; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_294;
  reg [7:0] _T_16959_37; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_295;
  reg [7:0] _T_16959_38; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_296;
  reg [7:0] _T_16959_39; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_297;
  reg [7:0] _T_16959_40; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_298;
  reg [7:0] _T_16959_41; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_299;
  reg [7:0] _T_16959_42; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_300;
  reg [7:0] _T_16959_43; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_301;
  reg [7:0] _T_16959_44; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_302;
  reg [7:0] _T_16959_45; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_303;
  reg [7:0] _T_16959_46; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_304;
  reg [7:0] _T_16959_47; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_305;
  reg [7:0] _T_16959_48; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_306;
  reg [7:0] _T_16959_49; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_307;
  reg [7:0] _T_16959_50; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_308;
  reg [7:0] _T_16959_51; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_309;
  reg [7:0] _T_16959_52; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_310;
  reg [7:0] _T_16959_53; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_311;
  reg [7:0] _T_16959_54; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_312;
  reg [7:0] _T_16959_55; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_313;
  reg [7:0] _T_16959_56; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_314;
  reg [7:0] _T_16959_57; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_315;
  reg [7:0] _T_16959_58; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_316;
  reg [7:0] _T_16959_59; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_317;
  reg [7:0] _T_16959_60; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_318;
  reg [7:0] _T_16959_61; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_319;
  reg [7:0] _T_16959_62; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_320;
  reg [7:0] _T_16959_63; // @[NV_NVDLA_CSC_WL_dec.scala 121:26:@13565.4]
  reg [31:0] _RAND_321;
  wire  _GEN_224; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_225; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_226; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_227; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_228; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_229; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_230; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_231; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_232; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_233; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_234; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_235; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_236; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_237; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_238; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_239; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_240; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_241; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_242; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_243; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_244; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_245; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_246; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_247; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_248; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_249; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_250; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_251; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_252; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_253; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_254; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire  _GEN_255; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  wire [7:0] _GEN_256; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13602.6]
  wire [7:0] _GEN_258; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13610.6]
  wire [7:0] _GEN_260; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13618.6]
  wire [7:0] _GEN_262; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13626.6]
  wire [7:0] _GEN_264; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13634.6]
  wire [7:0] _GEN_266; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13642.6]
  wire [7:0] _GEN_268; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13650.6]
  wire [7:0] _GEN_270; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13658.6]
  wire [7:0] _GEN_272; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13666.6]
  wire [7:0] _GEN_274; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13674.6]
  wire [7:0] _GEN_276; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13682.6]
  wire [7:0] _GEN_278; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13690.6]
  wire [7:0] _GEN_280; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13698.6]
  wire [7:0] _GEN_282; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13706.6]
  wire [7:0] _GEN_284; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13714.6]
  wire [7:0] _GEN_286; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13722.6]
  wire [7:0] _GEN_288; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13730.6]
  wire [7:0] _GEN_290; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13738.6]
  wire [7:0] _GEN_292; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13746.6]
  wire [7:0] _GEN_294; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13754.6]
  wire [7:0] _GEN_296; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13762.6]
  wire [7:0] _GEN_298; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13770.6]
  wire [7:0] _GEN_300; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13778.6]
  wire [7:0] _GEN_302; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13786.6]
  wire [7:0] _GEN_304; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13794.6]
  wire [7:0] _GEN_306; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13802.6]
  wire [7:0] _GEN_308; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13810.6]
  wire [7:0] _GEN_310; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13818.6]
  wire [7:0] _GEN_312; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13826.6]
  wire [7:0] _GEN_314; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13834.6]
  wire [7:0] _GEN_316; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13842.6]
  wire [7:0] _GEN_318; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13850.6]
  wire [7:0] _GEN_320; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13858.6]
  wire [7:0] _GEN_322; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13866.6]
  wire [7:0] _GEN_324; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13874.6]
  wire [7:0] _GEN_326; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13882.6]
  wire [7:0] _GEN_328; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13890.6]
  wire [7:0] _GEN_330; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13898.6]
  wire [7:0] _GEN_332; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13906.6]
  wire [7:0] _GEN_334; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13914.6]
  wire [7:0] _GEN_336; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13922.6]
  wire [7:0] _GEN_338; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13930.6]
  wire [7:0] _GEN_340; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13938.6]
  wire [7:0] _GEN_342; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13946.6]
  wire [7:0] _GEN_344; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13954.6]
  wire [7:0] _GEN_346; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13962.6]
  wire [7:0] _GEN_348; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13970.6]
  wire [7:0] _GEN_350; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13978.6]
  wire [7:0] _GEN_352; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13986.6]
  wire [7:0] _GEN_354; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13994.6]
  wire [7:0] _GEN_356; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14002.6]
  wire [7:0] _GEN_358; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14010.6]
  wire [7:0] _GEN_360; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14018.6]
  wire [7:0] _GEN_362; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14026.6]
  wire [7:0] _GEN_364; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14034.6]
  wire [7:0] _GEN_366; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14042.6]
  wire [7:0] _GEN_368; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14050.6]
  wire [7:0] _GEN_370; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14058.6]
  wire [7:0] _GEN_372; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14066.6]
  wire [7:0] _GEN_374; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14074.6]
  wire [7:0] _GEN_376; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14082.6]
  wire [7:0] _GEN_378; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14090.6]
  wire [7:0] _GEN_380; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14098.6]
  wire [7:0] _GEN_382; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14106.6]
  wire  _T_17161; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14114.4]
  wire  _T_17163; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14116.4]
  wire  _T_17165; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14118.4]
  wire  _T_17167; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14120.4]
  wire  _T_17169; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14122.4]
  wire  _T_17171; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14124.4]
  wire  _T_17173; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14126.4]
  wire  _T_17175; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14128.4]
  wire  _T_17177; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14130.4]
  wire  _T_17179; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14132.4]
  wire  _T_17181; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14134.4]
  wire  _T_17183; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14136.4]
  wire  _T_17185; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14138.4]
  wire  _T_17187; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14140.4]
  wire  _T_17189; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14142.4]
  wire  _T_17191; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14144.4]
  wire  _T_17193; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14146.4]
  wire  _T_17195; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14148.4]
  wire  _T_17197; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14150.4]
  wire  _T_17199; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14152.4]
  wire  _T_17201; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14154.4]
  wire  _T_17203; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14156.4]
  wire  _T_17205; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14158.4]
  wire  _T_17207; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14160.4]
  wire  _T_17209; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14162.4]
  wire  _T_17211; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14164.4]
  wire  _T_17213; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14166.4]
  wire  _T_17215; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14168.4]
  wire  _T_17217; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14170.4]
  wire  _T_17219; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14172.4]
  wire  _T_17221; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14174.4]
  wire  _T_17223; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14176.4]
  wire  _T_17225; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14178.4]
  wire  _T_17227; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14180.4]
  wire  _T_17229; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14182.4]
  wire  _T_17231; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14184.4]
  wire  _T_17233; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14186.4]
  wire  _T_17235; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14188.4]
  wire  _T_17237; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14190.4]
  wire  _T_17239; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14192.4]
  wire  _T_17241; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14194.4]
  wire  _T_17243; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14196.4]
  wire  _T_17245; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14198.4]
  wire  _T_17247; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14200.4]
  wire  _T_17249; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14202.4]
  wire  _T_17251; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14204.4]
  wire  _T_17253; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14206.4]
  wire  _T_17255; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14208.4]
  wire  _T_17257; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14210.4]
  wire  _T_17259; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14212.4]
  wire  _T_17261; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14214.4]
  wire  _T_17263; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14216.4]
  wire  _T_17265; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14218.4]
  wire  _T_17267; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14220.4]
  wire  _T_17269; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14222.4]
  wire  _T_17271; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14224.4]
  wire  _T_17273; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14226.4]
  wire  _T_17275; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14228.4]
  wire  _T_17277; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14230.4]
  wire  _T_17279; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14232.4]
  wire  _T_17281; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14234.4]
  wire  _T_17283; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14236.4]
  wire  _T_17285; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14238.4]
  wire  _T_17287; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14240.4]
  reg  _T_17290; // @[NV_NVDLA_CSC_WL_dec.scala 147:27:@14242.4]
  reg [31:0] _RAND_322;
  reg  _T_17294_0; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_323;
  reg  _T_17294_1; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_324;
  reg  _T_17294_2; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_325;
  reg  _T_17294_3; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_326;
  reg  _T_17294_4; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_327;
  reg  _T_17294_5; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_328;
  reg  _T_17294_6; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_329;
  reg  _T_17294_7; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_330;
  reg  _T_17294_8; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_331;
  reg  _T_17294_9; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_332;
  reg  _T_17294_10; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_333;
  reg  _T_17294_11; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_334;
  reg  _T_17294_12; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_335;
  reg  _T_17294_13; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_336;
  reg  _T_17294_14; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_337;
  reg  _T_17294_15; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_338;
  reg  _T_17294_16; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_339;
  reg  _T_17294_17; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_340;
  reg  _T_17294_18; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_341;
  reg  _T_17294_19; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_342;
  reg  _T_17294_20; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_343;
  reg  _T_17294_21; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_344;
  reg  _T_17294_22; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_345;
  reg  _T_17294_23; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_346;
  reg  _T_17294_24; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_347;
  reg  _T_17294_25; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_348;
  reg  _T_17294_26; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_349;
  reg  _T_17294_27; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_350;
  reg  _T_17294_28; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_351;
  reg  _T_17294_29; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_352;
  reg  _T_17294_30; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_353;
  reg  _T_17294_31; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_354;
  reg  _T_17294_32; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_355;
  reg  _T_17294_33; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_356;
  reg  _T_17294_34; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_357;
  reg  _T_17294_35; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_358;
  reg  _T_17294_36; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_359;
  reg  _T_17294_37; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_360;
  reg  _T_17294_38; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_361;
  reg  _T_17294_39; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_362;
  reg  _T_17294_40; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_363;
  reg  _T_17294_41; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_364;
  reg  _T_17294_42; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_365;
  reg  _T_17294_43; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_366;
  reg  _T_17294_44; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_367;
  reg  _T_17294_45; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_368;
  reg  _T_17294_46; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_369;
  reg  _T_17294_47; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_370;
  reg  _T_17294_48; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_371;
  reg  _T_17294_49; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_372;
  reg  _T_17294_50; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_373;
  reg  _T_17294_51; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_374;
  reg  _T_17294_52; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_375;
  reg  _T_17294_53; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_376;
  reg  _T_17294_54; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_377;
  reg  _T_17294_55; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_378;
  reg  _T_17294_56; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_379;
  reg  _T_17294_57; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_380;
  reg  _T_17294_58; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_381;
  reg  _T_17294_59; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_382;
  reg  _T_17294_60; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_383;
  reg  _T_17294_61; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_384;
  reg  _T_17294_62; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_385;
  reg  _T_17294_63; // @[NV_NVDLA_CSC_WL_dec.scala 148:22:@14243.4]
  reg [31:0] _RAND_386;
  reg  _T_17499_0; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_387;
  reg  _T_17499_1; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_388;
  reg  _T_17499_2; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_389;
  reg  _T_17499_3; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_390;
  reg  _T_17499_4; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_391;
  reg  _T_17499_5; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_392;
  reg  _T_17499_6; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_393;
  reg  _T_17499_7; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_394;
  reg  _T_17499_8; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_395;
  reg  _T_17499_9; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_396;
  reg  _T_17499_10; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_397;
  reg  _T_17499_11; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_398;
  reg  _T_17499_12; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_399;
  reg  _T_17499_13; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_400;
  reg  _T_17499_14; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_401;
  reg  _T_17499_15; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_402;
  reg  _T_17499_16; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_403;
  reg  _T_17499_17; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_404;
  reg  _T_17499_18; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_405;
  reg  _T_17499_19; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_406;
  reg  _T_17499_20; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_407;
  reg  _T_17499_21; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_408;
  reg  _T_17499_22; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_409;
  reg  _T_17499_23; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_410;
  reg  _T_17499_24; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_411;
  reg  _T_17499_25; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_412;
  reg  _T_17499_26; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_413;
  reg  _T_17499_27; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_414;
  reg  _T_17499_28; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_415;
  reg  _T_17499_29; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_416;
  reg  _T_17499_30; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_417;
  reg  _T_17499_31; // @[NV_NVDLA_CSC_WL_dec.scala 149:25:@14277.4]
  reg [31:0] _RAND_418;
  reg [7:0] _T_17603_0; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_419;
  reg [7:0] _T_17603_1; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_420;
  reg [7:0] _T_17603_2; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_421;
  reg [7:0] _T_17603_3; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_422;
  reg [7:0] _T_17603_4; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_423;
  reg [7:0] _T_17603_5; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_424;
  reg [7:0] _T_17603_6; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_425;
  reg [7:0] _T_17603_7; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_426;
  reg [7:0] _T_17603_8; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_427;
  reg [7:0] _T_17603_9; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_428;
  reg [7:0] _T_17603_10; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_429;
  reg [7:0] _T_17603_11; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_430;
  reg [7:0] _T_17603_12; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_431;
  reg [7:0] _T_17603_13; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_432;
  reg [7:0] _T_17603_14; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_433;
  reg [7:0] _T_17603_15; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_434;
  reg [7:0] _T_17603_16; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_435;
  reg [7:0] _T_17603_17; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_436;
  reg [7:0] _T_17603_18; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_437;
  reg [7:0] _T_17603_19; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_438;
  reg [7:0] _T_17603_20; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_439;
  reg [7:0] _T_17603_21; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_440;
  reg [7:0] _T_17603_22; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_441;
  reg [7:0] _T_17603_23; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_442;
  reg [7:0] _T_17603_24; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_443;
  reg [7:0] _T_17603_25; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_444;
  reg [7:0] _T_17603_26; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_445;
  reg [7:0] _T_17603_27; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_446;
  reg [7:0] _T_17603_28; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_447;
  reg [7:0] _T_17603_29; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_448;
  reg [7:0] _T_17603_30; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_449;
  reg [7:0] _T_17603_31; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_450;
  reg [7:0] _T_17603_32; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_451;
  reg [7:0] _T_17603_33; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_452;
  reg [7:0] _T_17603_34; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_453;
  reg [7:0] _T_17603_35; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_454;
  reg [7:0] _T_17603_36; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_455;
  reg [7:0] _T_17603_37; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_456;
  reg [7:0] _T_17603_38; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_457;
  reg [7:0] _T_17603_39; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_458;
  reg [7:0] _T_17603_40; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_459;
  reg [7:0] _T_17603_41; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_460;
  reg [7:0] _T_17603_42; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_461;
  reg [7:0] _T_17603_43; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_462;
  reg [7:0] _T_17603_44; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_463;
  reg [7:0] _T_17603_45; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_464;
  reg [7:0] _T_17603_46; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_465;
  reg [7:0] _T_17603_47; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_466;
  reg [7:0] _T_17603_48; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_467;
  reg [7:0] _T_17603_49; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_468;
  reg [7:0] _T_17603_50; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_469;
  reg [7:0] _T_17603_51; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_470;
  reg [7:0] _T_17603_52; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_471;
  reg [7:0] _T_17603_53; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_472;
  reg [7:0] _T_17603_54; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_473;
  reg [7:0] _T_17603_55; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_474;
  reg [7:0] _T_17603_56; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_475;
  reg [7:0] _T_17603_57; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_476;
  reg [7:0] _T_17603_58; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_477;
  reg [7:0] _T_17603_59; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_478;
  reg [7:0] _T_17603_60; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_479;
  reg [7:0] _T_17603_61; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_480;
  reg [7:0] _T_17603_62; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_481;
  reg [7:0] _T_17603_63; // @[NV_NVDLA_CSC_WL_dec.scala 150:26:@14278.4]
  reg [31:0] _RAND_482;
  wire  _GEN_448; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_449; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_450; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_451; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_452; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_453; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_454; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_455; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_456; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_457; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_458; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_459; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_460; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_461; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_462; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_463; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_464; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_465; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_466; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_467; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_468; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_469; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_470; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_471; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_472; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_473; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_474; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_475; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_476; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_477; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_478; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire  _GEN_479; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  wire [7:0] _T_17676; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14449.4]
  wire [15:0] _T_17684; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14457.4]
  wire [7:0] _T_17691; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14464.4]
  wire [31:0] _T_17700; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14473.4]
  wire [7:0] _T_17707; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14480.4]
  wire [15:0] _T_17715; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14488.4]
  wire [7:0] _T_17722; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14495.4]
  wire [31:0] _T_17731; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14504.4]
  wire [7:0] _T_17739; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14513.4]
  wire [15:0] _T_17747; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14521.4]
  wire [7:0] _T_17754; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14528.4]
  wire [15:0] _T_17762; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14536.4]
  assign _T_326 = io_nvdla_core_rstn == 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 55:37:@8.4]
  assign _T_397 = io_input_bits_mask[0]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@10.4]
  assign _T_398 = io_input_bits_mask[1]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@12.4]
  assign _T_399 = io_input_bits_mask[2]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@14.4]
  assign _T_400 = io_input_bits_mask[3]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@16.4]
  assign _T_401 = io_input_bits_mask[4]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@18.4]
  assign _T_402 = io_input_bits_mask[5]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@20.4]
  assign _T_403 = io_input_bits_mask[6]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@22.4]
  assign _T_404 = io_input_bits_mask[7]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@24.4]
  assign _T_405 = io_input_bits_mask[8]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@26.4]
  assign _T_406 = io_input_bits_mask[9]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@28.4]
  assign _T_407 = io_input_bits_mask[10]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@30.4]
  assign _T_408 = io_input_bits_mask[11]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@32.4]
  assign _T_409 = io_input_bits_mask[12]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@34.4]
  assign _T_410 = io_input_bits_mask[13]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@36.4]
  assign _T_411 = io_input_bits_mask[14]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@38.4]
  assign _T_412 = io_input_bits_mask[15]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@40.4]
  assign _T_413 = io_input_bits_mask[16]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@42.4]
  assign _T_414 = io_input_bits_mask[17]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@44.4]
  assign _T_415 = io_input_bits_mask[18]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@46.4]
  assign _T_416 = io_input_bits_mask[19]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@48.4]
  assign _T_417 = io_input_bits_mask[20]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@50.4]
  assign _T_418 = io_input_bits_mask[21]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@52.4]
  assign _T_419 = io_input_bits_mask[22]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@54.4]
  assign _T_420 = io_input_bits_mask[23]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@56.4]
  assign _T_421 = io_input_bits_mask[24]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@58.4]
  assign _T_422 = io_input_bits_mask[25]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@60.4]
  assign _T_423 = io_input_bits_mask[26]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@62.4]
  assign _T_424 = io_input_bits_mask[27]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@64.4]
  assign _T_425 = io_input_bits_mask[28]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@66.4]
  assign _T_426 = io_input_bits_mask[29]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@68.4]
  assign _T_427 = io_input_bits_mask[30]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@70.4]
  assign _T_428 = io_input_bits_mask[31]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@72.4]
  assign _T_429 = io_input_bits_mask[32]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@74.4]
  assign _T_430 = io_input_bits_mask[33]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@76.4]
  assign _T_431 = io_input_bits_mask[34]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@78.4]
  assign _T_432 = io_input_bits_mask[35]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@80.4]
  assign _T_433 = io_input_bits_mask[36]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@82.4]
  assign _T_434 = io_input_bits_mask[37]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@84.4]
  assign _T_435 = io_input_bits_mask[38]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@86.4]
  assign _T_436 = io_input_bits_mask[39]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@88.4]
  assign _T_437 = io_input_bits_mask[40]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@90.4]
  assign _T_438 = io_input_bits_mask[41]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@92.4]
  assign _T_439 = io_input_bits_mask[42]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@94.4]
  assign _T_440 = io_input_bits_mask[43]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@96.4]
  assign _T_441 = io_input_bits_mask[44]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@98.4]
  assign _T_442 = io_input_bits_mask[45]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@100.4]
  assign _T_443 = io_input_bits_mask[46]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@102.4]
  assign _T_444 = io_input_bits_mask[47]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@104.4]
  assign _T_445 = io_input_bits_mask[48]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@106.4]
  assign _T_446 = io_input_bits_mask[49]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@108.4]
  assign _T_447 = io_input_bits_mask[50]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@110.4]
  assign _T_448 = io_input_bits_mask[51]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@112.4]
  assign _T_449 = io_input_bits_mask[52]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@114.4]
  assign _T_450 = io_input_bits_mask[53]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@116.4]
  assign _T_451 = io_input_bits_mask[54]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@118.4]
  assign _T_452 = io_input_bits_mask[55]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@120.4]
  assign _T_453 = io_input_bits_mask[56]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@122.4]
  assign _T_454 = io_input_bits_mask[57]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@124.4]
  assign _T_455 = io_input_bits_mask[58]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@126.4]
  assign _T_456 = io_input_bits_mask[59]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@128.4]
  assign _T_457 = io_input_bits_mask[60]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@130.4]
  assign _T_458 = io_input_bits_mask[61]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@132.4]
  assign _T_459 = io_input_bits_mask[62]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@134.4]
  assign _T_460 = io_input_bits_mask[63]; // @[NV_NVDLA_CSC_WL_dec.scala 70:48:@136.4]
  assign _T_531 = io_input_bits_data[7:0]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@139.4]
  assign _T_532 = io_input_bits_data[15:8]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@141.4]
  assign _T_533 = io_input_bits_data[23:16]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@143.4]
  assign _T_534 = io_input_bits_data[31:24]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@145.4]
  assign _T_535 = io_input_bits_data[39:32]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@147.4]
  assign _T_536 = io_input_bits_data[47:40]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@149.4]
  assign _T_537 = io_input_bits_data[55:48]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@151.4]
  assign _T_538 = io_input_bits_data[63:56]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@153.4]
  assign _T_539 = io_input_bits_data[71:64]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@155.4]
  assign _T_540 = io_input_bits_data[79:72]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@157.4]
  assign _T_541 = io_input_bits_data[87:80]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@159.4]
  assign _T_542 = io_input_bits_data[95:88]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@161.4]
  assign _T_543 = io_input_bits_data[103:96]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@163.4]
  assign _T_544 = io_input_bits_data[111:104]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@165.4]
  assign _T_545 = io_input_bits_data[119:112]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@167.4]
  assign _T_546 = io_input_bits_data[127:120]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@169.4]
  assign _T_547 = io_input_bits_data[135:128]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@171.4]
  assign _T_548 = io_input_bits_data[143:136]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@173.4]
  assign _T_549 = io_input_bits_data[151:144]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@175.4]
  assign _T_550 = io_input_bits_data[159:152]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@177.4]
  assign _T_551 = io_input_bits_data[167:160]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@179.4]
  assign _T_552 = io_input_bits_data[175:168]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@181.4]
  assign _T_553 = io_input_bits_data[183:176]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@183.4]
  assign _T_554 = io_input_bits_data[191:184]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@185.4]
  assign _T_555 = io_input_bits_data[199:192]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@187.4]
  assign _T_556 = io_input_bits_data[207:200]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@189.4]
  assign _T_557 = io_input_bits_data[215:208]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@191.4]
  assign _T_558 = io_input_bits_data[223:216]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@193.4]
  assign _T_559 = io_input_bits_data[231:224]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@195.4]
  assign _T_560 = io_input_bits_data[239:232]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@197.4]
  assign _T_561 = io_input_bits_data[247:240]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@199.4]
  assign _T_562 = io_input_bits_data[255:248]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@201.4]
  assign _T_563 = io_input_bits_data[263:256]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@203.4]
  assign _T_564 = io_input_bits_data[271:264]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@205.4]
  assign _T_565 = io_input_bits_data[279:272]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@207.4]
  assign _T_566 = io_input_bits_data[287:280]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@209.4]
  assign _T_567 = io_input_bits_data[295:288]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@211.4]
  assign _T_568 = io_input_bits_data[303:296]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@213.4]
  assign _T_569 = io_input_bits_data[311:304]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@215.4]
  assign _T_570 = io_input_bits_data[319:312]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@217.4]
  assign _T_571 = io_input_bits_data[327:320]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@219.4]
  assign _T_572 = io_input_bits_data[335:328]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@221.4]
  assign _T_573 = io_input_bits_data[343:336]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@223.4]
  assign _T_574 = io_input_bits_data[351:344]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@225.4]
  assign _T_575 = io_input_bits_data[359:352]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@227.4]
  assign _T_576 = io_input_bits_data[367:360]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@229.4]
  assign _T_577 = io_input_bits_data[375:368]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@231.4]
  assign _T_578 = io_input_bits_data[383:376]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@233.4]
  assign _T_579 = io_input_bits_data[391:384]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@235.4]
  assign _T_580 = io_input_bits_data[399:392]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@237.4]
  assign _T_581 = io_input_bits_data[407:400]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@239.4]
  assign _T_582 = io_input_bits_data[415:408]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@241.4]
  assign _T_583 = io_input_bits_data[423:416]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@243.4]
  assign _T_584 = io_input_bits_data[431:424]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@245.4]
  assign _T_585 = io_input_bits_data[439:432]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@247.4]
  assign _T_586 = io_input_bits_data[447:440]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@249.4]
  assign _T_587 = io_input_bits_data[455:448]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@251.4]
  assign _T_588 = io_input_bits_data[463:456]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@253.4]
  assign _T_589 = io_input_bits_data[471:464]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@255.4]
  assign _T_590 = io_input_bits_data[479:472]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@257.4]
  assign _T_591 = io_input_bits_data[487:480]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@259.4]
  assign _T_592 = io_input_bits_data[495:488]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@261.4]
  assign _T_593 = io_input_bits_data[503:496]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@263.4]
  assign _T_594 = io_input_bits_data[511:504]; // @[NV_NVDLA_CSC_WL_dec.scala 74:48:@265.4]
  assign _T_633 = io_input_bits_sel[0]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@268.4]
  assign _T_634 = io_input_bits_sel[1]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@270.4]
  assign _T_635 = io_input_bits_sel[2]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@272.4]
  assign _T_636 = io_input_bits_sel[3]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@274.4]
  assign _T_637 = io_input_bits_sel[4]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@276.4]
  assign _T_638 = io_input_bits_sel[5]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@278.4]
  assign _T_639 = io_input_bits_sel[6]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@280.4]
  assign _T_640 = io_input_bits_sel[7]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@282.4]
  assign _T_641 = io_input_bits_sel[8]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@284.4]
  assign _T_642 = io_input_bits_sel[9]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@286.4]
  assign _T_643 = io_input_bits_sel[10]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@288.4]
  assign _T_644 = io_input_bits_sel[11]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@290.4]
  assign _T_645 = io_input_bits_sel[12]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@292.4]
  assign _T_646 = io_input_bits_sel[13]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@294.4]
  assign _T_647 = io_input_bits_sel[14]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@296.4]
  assign _T_648 = io_input_bits_sel[15]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@298.4]
  assign _T_649 = io_input_bits_sel[16]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@300.4]
  assign _T_650 = io_input_bits_sel[17]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@302.4]
  assign _T_651 = io_input_bits_sel[18]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@304.4]
  assign _T_652 = io_input_bits_sel[19]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@306.4]
  assign _T_653 = io_input_bits_sel[20]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@308.4]
  assign _T_654 = io_input_bits_sel[21]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@310.4]
  assign _T_655 = io_input_bits_sel[22]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@312.4]
  assign _T_656 = io_input_bits_sel[23]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@314.4]
  assign _T_657 = io_input_bits_sel[24]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@316.4]
  assign _T_658 = io_input_bits_sel[25]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@318.4]
  assign _T_659 = io_input_bits_sel[26]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@320.4]
  assign _T_660 = io_input_bits_sel[27]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@322.4]
  assign _T_661 = io_input_bits_sel[28]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@324.4]
  assign _T_662 = io_input_bits_sel[29]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@326.4]
  assign _T_663 = io_input_bits_sel[30]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@328.4]
  assign _T_664 = io_input_bits_sel[31]; // @[NV_NVDLA_CSC_WL_dec.scala 78:46:@330.4]
  assign _T_665 = io_input_mask_en[8]; // @[NV_NVDLA_CSC_WL_dec.scala 81:48:@332.4]
  assign _T_800_0 = _T_665 ? _T_397 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_1 = _T_665 ? _T_398 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_2 = _T_665 ? _T_399 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_3 = _T_665 ? _T_400 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_4 = _T_665 ? _T_401 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_5 = _T_665 ? _T_402 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_6 = _T_665 ? _T_403 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_7 = _T_665 ? _T_404 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_8 = _T_665 ? _T_405 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_9 = _T_665 ? _T_406 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_10 = _T_665 ? _T_407 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_11 = _T_665 ? _T_408 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_12 = _T_665 ? _T_409 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_13 = _T_665 ? _T_410 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_14 = _T_665 ? _T_411 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_15 = _T_665 ? _T_412 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_16 = _T_665 ? _T_413 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_17 = _T_665 ? _T_414 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_18 = _T_665 ? _T_415 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_19 = _T_665 ? _T_416 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_20 = _T_665 ? _T_417 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_21 = _T_665 ? _T_418 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_22 = _T_665 ? _T_419 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_23 = _T_665 ? _T_420 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_24 = _T_665 ? _T_421 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_25 = _T_665 ? _T_422 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_26 = _T_665 ? _T_423 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_27 = _T_665 ? _T_424 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_28 = _T_665 ? _T_425 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_29 = _T_665 ? _T_426 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_30 = _T_665 ? _T_427 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_31 = _T_665 ? _T_428 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_32 = _T_665 ? _T_429 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_33 = _T_665 ? _T_430 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_34 = _T_665 ? _T_431 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_35 = _T_665 ? _T_432 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_36 = _T_665 ? _T_433 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_37 = _T_665 ? _T_434 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_38 = _T_665 ? _T_435 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_39 = _T_665 ? _T_436 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_40 = _T_665 ? _T_437 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_41 = _T_665 ? _T_438 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_42 = _T_665 ? _T_439 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_43 = _T_665 ? _T_440 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_44 = _T_665 ? _T_441 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_45 = _T_665 ? _T_442 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_46 = _T_665 ? _T_443 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_47 = _T_665 ? _T_444 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_48 = _T_665 ? _T_445 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_49 = _T_665 ? _T_446 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_50 = _T_665 ? _T_447 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_51 = _T_665 ? _T_448 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_52 = _T_665 ? _T_449 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_53 = _T_665 ? _T_450 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_54 = _T_665 ? _T_451 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_55 = _T_665 ? _T_452 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_56 = _T_665 ? _T_453 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_57 = _T_665 ? _T_454 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_58 = _T_665 ? _T_455 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_59 = _T_665 ? _T_456 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_60 = _T_665 ? _T_457 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_61 = _T_665 ? _T_458 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_62 = _T_665 ? _T_459 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_800_63 = _T_665 ? _T_460 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 81:31:@398.4]
  assign _T_1068 = {_T_800_7,_T_800_6,_T_800_5,_T_800_4,_T_800_3,_T_800_2,_T_800_1,_T_800_0}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@406.4]
  assign _T_1076 = {_T_800_15,_T_800_14,_T_800_13,_T_800_12,_T_800_11,_T_800_10,_T_800_9,_T_800_8,_T_1068}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@414.4]
  assign _T_1083 = {_T_800_23,_T_800_22,_T_800_21,_T_800_20,_T_800_19,_T_800_18,_T_800_17,_T_800_16}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@421.4]
  assign _T_1092 = {_T_800_31,_T_800_30,_T_800_29,_T_800_28,_T_800_27,_T_800_26,_T_800_25,_T_800_24,_T_1083,_T_1076}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@430.4]
  assign _T_1099 = {_T_800_39,_T_800_38,_T_800_37,_T_800_36,_T_800_35,_T_800_34,_T_800_33,_T_800_32}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@437.4]
  assign _T_1107 = {_T_800_47,_T_800_46,_T_800_45,_T_800_44,_T_800_43,_T_800_42,_T_800_41,_T_800_40,_T_1099}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@445.4]
  assign _T_1114 = {_T_800_55,_T_800_54,_T_800_53,_T_800_52,_T_800_51,_T_800_50,_T_800_49,_T_800_48}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@452.4]
  assign _T_1123 = {_T_800_63,_T_800_62,_T_800_61,_T_800_60,_T_800_59,_T_800_58,_T_800_57,_T_800_56,_T_1114,_T_1107}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@461.4]
  assign _T_1124 = {_T_1123,_T_1092}; // @[NV_NVDLA_CSC_WL_dec.scala 85:53:@462.4]
  assign _T_1125 = _T_1124[0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@463.4]
  assign _T_1190 = _T_1124[1:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@529.4]
  assign _T_1191 = _T_1190[0]; // @[Bitwise.scala 50:65:@530.4]
  assign _T_1192 = _T_1190[1]; // @[Bitwise.scala 50:65:@531.4]
  assign _T_1193 = _T_1191 + _T_1192; // @[Bitwise.scala 48:55:@532.4]
  assign _T_1257 = _T_1124[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@597.4]
  assign _T_1258 = _T_1257[0]; // @[Bitwise.scala 50:65:@598.4]
  assign _T_1259 = _T_1257[1]; // @[Bitwise.scala 50:65:@599.4]
  assign _T_1260 = _T_1257[2]; // @[Bitwise.scala 50:65:@600.4]
  assign _T_1261 = _T_1259 + _T_1260; // @[Bitwise.scala 48:55:@601.4]
  assign _GEN_544 = {{1'd0}, _T_1258}; // @[Bitwise.scala 48:55:@602.4]
  assign _T_1262 = _GEN_544 + _T_1261; // @[Bitwise.scala 48:55:@602.4]
  assign _T_1326 = _T_1124[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@667.4]
  assign _T_1327 = _T_1326[0]; // @[Bitwise.scala 50:65:@668.4]
  assign _T_1328 = _T_1326[1]; // @[Bitwise.scala 50:65:@669.4]
  assign _T_1329 = _T_1326[2]; // @[Bitwise.scala 50:65:@670.4]
  assign _T_1330 = _T_1326[3]; // @[Bitwise.scala 50:65:@671.4]
  assign _T_1331 = _T_1327 + _T_1328; // @[Bitwise.scala 48:55:@672.4]
  assign _T_1332 = _T_1329 + _T_1330; // @[Bitwise.scala 48:55:@673.4]
  assign _T_1333 = _T_1331 + _T_1332; // @[Bitwise.scala 48:55:@674.4]
  assign _T_1397 = _T_1124[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@739.4]
  assign _T_1398 = _T_1397[0]; // @[Bitwise.scala 50:65:@740.4]
  assign _T_1399 = _T_1397[1]; // @[Bitwise.scala 50:65:@741.4]
  assign _T_1400 = _T_1397[2]; // @[Bitwise.scala 50:65:@742.4]
  assign _T_1401 = _T_1397[3]; // @[Bitwise.scala 50:65:@743.4]
  assign _T_1402 = _T_1397[4]; // @[Bitwise.scala 50:65:@744.4]
  assign _T_1403 = _T_1398 + _T_1399; // @[Bitwise.scala 48:55:@745.4]
  assign _T_1404 = _T_1401 + _T_1402; // @[Bitwise.scala 48:55:@746.4]
  assign _GEN_545 = {{1'd0}, _T_1400}; // @[Bitwise.scala 48:55:@747.4]
  assign _T_1405 = _GEN_545 + _T_1404; // @[Bitwise.scala 48:55:@747.4]
  assign _GEN_546 = {{1'd0}, _T_1403}; // @[Bitwise.scala 48:55:@748.4]
  assign _T_1406 = _GEN_546 + _T_1405; // @[Bitwise.scala 48:55:@748.4]
  assign _T_1470 = _T_1124[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@813.4]
  assign _T_1471 = _T_1470[0]; // @[Bitwise.scala 50:65:@814.4]
  assign _T_1472 = _T_1470[1]; // @[Bitwise.scala 50:65:@815.4]
  assign _T_1473 = _T_1470[2]; // @[Bitwise.scala 50:65:@816.4]
  assign _T_1474 = _T_1470[3]; // @[Bitwise.scala 50:65:@817.4]
  assign _T_1475 = _T_1470[4]; // @[Bitwise.scala 50:65:@818.4]
  assign _T_1476 = _T_1470[5]; // @[Bitwise.scala 50:65:@819.4]
  assign _T_1477 = _T_1472 + _T_1473; // @[Bitwise.scala 48:55:@820.4]
  assign _GEN_547 = {{1'd0}, _T_1471}; // @[Bitwise.scala 48:55:@821.4]
  assign _T_1478 = _GEN_547 + _T_1477; // @[Bitwise.scala 48:55:@821.4]
  assign _T_1479 = _T_1475 + _T_1476; // @[Bitwise.scala 48:55:@822.4]
  assign _GEN_548 = {{1'd0}, _T_1474}; // @[Bitwise.scala 48:55:@823.4]
  assign _T_1480 = _GEN_548 + _T_1479; // @[Bitwise.scala 48:55:@823.4]
  assign _T_1481 = _T_1478 + _T_1480; // @[Bitwise.scala 48:55:@824.4]
  assign _T_1545 = _T_1124[6:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@889.4]
  assign _T_1546 = _T_1545[0]; // @[Bitwise.scala 50:65:@890.4]
  assign _T_1547 = _T_1545[1]; // @[Bitwise.scala 50:65:@891.4]
  assign _T_1548 = _T_1545[2]; // @[Bitwise.scala 50:65:@892.4]
  assign _T_1549 = _T_1545[3]; // @[Bitwise.scala 50:65:@893.4]
  assign _T_1550 = _T_1545[4]; // @[Bitwise.scala 50:65:@894.4]
  assign _T_1551 = _T_1545[5]; // @[Bitwise.scala 50:65:@895.4]
  assign _T_1552 = _T_1545[6]; // @[Bitwise.scala 50:65:@896.4]
  assign _T_1553 = _T_1547 + _T_1548; // @[Bitwise.scala 48:55:@897.4]
  assign _GEN_549 = {{1'd0}, _T_1546}; // @[Bitwise.scala 48:55:@898.4]
  assign _T_1554 = _GEN_549 + _T_1553; // @[Bitwise.scala 48:55:@898.4]
  assign _T_1555 = _T_1549 + _T_1550; // @[Bitwise.scala 48:55:@899.4]
  assign _T_1556 = _T_1551 + _T_1552; // @[Bitwise.scala 48:55:@900.4]
  assign _T_1557 = _T_1555 + _T_1556; // @[Bitwise.scala 48:55:@901.4]
  assign _T_1558 = _T_1554 + _T_1557; // @[Bitwise.scala 48:55:@902.4]
  assign _T_1622 = _T_1124[7:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@967.4]
  assign _T_1623 = _T_1622[0]; // @[Bitwise.scala 50:65:@968.4]
  assign _T_1624 = _T_1622[1]; // @[Bitwise.scala 50:65:@969.4]
  assign _T_1625 = _T_1622[2]; // @[Bitwise.scala 50:65:@970.4]
  assign _T_1626 = _T_1622[3]; // @[Bitwise.scala 50:65:@971.4]
  assign _T_1627 = _T_1622[4]; // @[Bitwise.scala 50:65:@972.4]
  assign _T_1628 = _T_1622[5]; // @[Bitwise.scala 50:65:@973.4]
  assign _T_1629 = _T_1622[6]; // @[Bitwise.scala 50:65:@974.4]
  assign _T_1630 = _T_1622[7]; // @[Bitwise.scala 50:65:@975.4]
  assign _T_1631 = _T_1623 + _T_1624; // @[Bitwise.scala 48:55:@976.4]
  assign _T_1632 = _T_1625 + _T_1626; // @[Bitwise.scala 48:55:@977.4]
  assign _T_1633 = _T_1631 + _T_1632; // @[Bitwise.scala 48:55:@978.4]
  assign _T_1634 = _T_1627 + _T_1628; // @[Bitwise.scala 48:55:@979.4]
  assign _T_1635 = _T_1629 + _T_1630; // @[Bitwise.scala 48:55:@980.4]
  assign _T_1636 = _T_1634 + _T_1635; // @[Bitwise.scala 48:55:@981.4]
  assign _T_1637 = _T_1633 + _T_1636; // @[Bitwise.scala 48:55:@982.4]
  assign _T_1701 = _T_1124[8:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1047.4]
  assign _T_1702 = _T_1701[0]; // @[Bitwise.scala 50:65:@1048.4]
  assign _T_1703 = _T_1701[1]; // @[Bitwise.scala 50:65:@1049.4]
  assign _T_1704 = _T_1701[2]; // @[Bitwise.scala 50:65:@1050.4]
  assign _T_1705 = _T_1701[3]; // @[Bitwise.scala 50:65:@1051.4]
  assign _T_1706 = _T_1701[4]; // @[Bitwise.scala 50:65:@1052.4]
  assign _T_1707 = _T_1701[5]; // @[Bitwise.scala 50:65:@1053.4]
  assign _T_1708 = _T_1701[6]; // @[Bitwise.scala 50:65:@1054.4]
  assign _T_1709 = _T_1701[7]; // @[Bitwise.scala 50:65:@1055.4]
  assign _T_1710 = _T_1701[8]; // @[Bitwise.scala 50:65:@1056.4]
  assign _T_1711 = _T_1702 + _T_1703; // @[Bitwise.scala 48:55:@1057.4]
  assign _T_1712 = _T_1704 + _T_1705; // @[Bitwise.scala 48:55:@1058.4]
  assign _T_1713 = _T_1711 + _T_1712; // @[Bitwise.scala 48:55:@1059.4]
  assign _T_1714 = _T_1706 + _T_1707; // @[Bitwise.scala 48:55:@1060.4]
  assign _T_1715 = _T_1709 + _T_1710; // @[Bitwise.scala 48:55:@1061.4]
  assign _GEN_550 = {{1'd0}, _T_1708}; // @[Bitwise.scala 48:55:@1062.4]
  assign _T_1716 = _GEN_550 + _T_1715; // @[Bitwise.scala 48:55:@1062.4]
  assign _GEN_551 = {{1'd0}, _T_1714}; // @[Bitwise.scala 48:55:@1063.4]
  assign _T_1717 = _GEN_551 + _T_1716; // @[Bitwise.scala 48:55:@1063.4]
  assign _GEN_552 = {{1'd0}, _T_1713}; // @[Bitwise.scala 48:55:@1064.4]
  assign _T_1718 = _GEN_552 + _T_1717; // @[Bitwise.scala 48:55:@1064.4]
  assign _T_1782 = _T_1124[9:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1129.4]
  assign _T_1783 = _T_1782[0]; // @[Bitwise.scala 50:65:@1130.4]
  assign _T_1784 = _T_1782[1]; // @[Bitwise.scala 50:65:@1131.4]
  assign _T_1785 = _T_1782[2]; // @[Bitwise.scala 50:65:@1132.4]
  assign _T_1786 = _T_1782[3]; // @[Bitwise.scala 50:65:@1133.4]
  assign _T_1787 = _T_1782[4]; // @[Bitwise.scala 50:65:@1134.4]
  assign _T_1788 = _T_1782[5]; // @[Bitwise.scala 50:65:@1135.4]
  assign _T_1789 = _T_1782[6]; // @[Bitwise.scala 50:65:@1136.4]
  assign _T_1790 = _T_1782[7]; // @[Bitwise.scala 50:65:@1137.4]
  assign _T_1791 = _T_1782[8]; // @[Bitwise.scala 50:65:@1138.4]
  assign _T_1792 = _T_1782[9]; // @[Bitwise.scala 50:65:@1139.4]
  assign _T_1793 = _T_1783 + _T_1784; // @[Bitwise.scala 48:55:@1140.4]
  assign _T_1794 = _T_1786 + _T_1787; // @[Bitwise.scala 48:55:@1141.4]
  assign _GEN_553 = {{1'd0}, _T_1785}; // @[Bitwise.scala 48:55:@1142.4]
  assign _T_1795 = _GEN_553 + _T_1794; // @[Bitwise.scala 48:55:@1142.4]
  assign _GEN_554 = {{1'd0}, _T_1793}; // @[Bitwise.scala 48:55:@1143.4]
  assign _T_1796 = _GEN_554 + _T_1795; // @[Bitwise.scala 48:55:@1143.4]
  assign _T_1797 = _T_1788 + _T_1789; // @[Bitwise.scala 48:55:@1144.4]
  assign _T_1798 = _T_1791 + _T_1792; // @[Bitwise.scala 48:55:@1145.4]
  assign _GEN_555 = {{1'd0}, _T_1790}; // @[Bitwise.scala 48:55:@1146.4]
  assign _T_1799 = _GEN_555 + _T_1798; // @[Bitwise.scala 48:55:@1146.4]
  assign _GEN_556 = {{1'd0}, _T_1797}; // @[Bitwise.scala 48:55:@1147.4]
  assign _T_1800 = _GEN_556 + _T_1799; // @[Bitwise.scala 48:55:@1147.4]
  assign _T_1801 = _T_1796 + _T_1800; // @[Bitwise.scala 48:55:@1148.4]
  assign _T_1865 = _T_1124[10:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1213.4]
  assign _T_1866 = _T_1865[0]; // @[Bitwise.scala 50:65:@1214.4]
  assign _T_1867 = _T_1865[1]; // @[Bitwise.scala 50:65:@1215.4]
  assign _T_1868 = _T_1865[2]; // @[Bitwise.scala 50:65:@1216.4]
  assign _T_1869 = _T_1865[3]; // @[Bitwise.scala 50:65:@1217.4]
  assign _T_1870 = _T_1865[4]; // @[Bitwise.scala 50:65:@1218.4]
  assign _T_1871 = _T_1865[5]; // @[Bitwise.scala 50:65:@1219.4]
  assign _T_1872 = _T_1865[6]; // @[Bitwise.scala 50:65:@1220.4]
  assign _T_1873 = _T_1865[7]; // @[Bitwise.scala 50:65:@1221.4]
  assign _T_1874 = _T_1865[8]; // @[Bitwise.scala 50:65:@1222.4]
  assign _T_1875 = _T_1865[9]; // @[Bitwise.scala 50:65:@1223.4]
  assign _T_1876 = _T_1865[10]; // @[Bitwise.scala 50:65:@1224.4]
  assign _T_1877 = _T_1866 + _T_1867; // @[Bitwise.scala 48:55:@1225.4]
  assign _T_1878 = _T_1869 + _T_1870; // @[Bitwise.scala 48:55:@1226.4]
  assign _GEN_557 = {{1'd0}, _T_1868}; // @[Bitwise.scala 48:55:@1227.4]
  assign _T_1879 = _GEN_557 + _T_1878; // @[Bitwise.scala 48:55:@1227.4]
  assign _GEN_558 = {{1'd0}, _T_1877}; // @[Bitwise.scala 48:55:@1228.4]
  assign _T_1880 = _GEN_558 + _T_1879; // @[Bitwise.scala 48:55:@1228.4]
  assign _T_1881 = _T_1872 + _T_1873; // @[Bitwise.scala 48:55:@1229.4]
  assign _GEN_559 = {{1'd0}, _T_1871}; // @[Bitwise.scala 48:55:@1230.4]
  assign _T_1882 = _GEN_559 + _T_1881; // @[Bitwise.scala 48:55:@1230.4]
  assign _T_1883 = _T_1875 + _T_1876; // @[Bitwise.scala 48:55:@1231.4]
  assign _GEN_560 = {{1'd0}, _T_1874}; // @[Bitwise.scala 48:55:@1232.4]
  assign _T_1884 = _GEN_560 + _T_1883; // @[Bitwise.scala 48:55:@1232.4]
  assign _T_1885 = _T_1882 + _T_1884; // @[Bitwise.scala 48:55:@1233.4]
  assign _T_1886 = _T_1880 + _T_1885; // @[Bitwise.scala 48:55:@1234.4]
  assign _T_1950 = _T_1124[11:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1299.4]
  assign _T_1951 = _T_1950[0]; // @[Bitwise.scala 50:65:@1300.4]
  assign _T_1952 = _T_1950[1]; // @[Bitwise.scala 50:65:@1301.4]
  assign _T_1953 = _T_1950[2]; // @[Bitwise.scala 50:65:@1302.4]
  assign _T_1954 = _T_1950[3]; // @[Bitwise.scala 50:65:@1303.4]
  assign _T_1955 = _T_1950[4]; // @[Bitwise.scala 50:65:@1304.4]
  assign _T_1956 = _T_1950[5]; // @[Bitwise.scala 50:65:@1305.4]
  assign _T_1957 = _T_1950[6]; // @[Bitwise.scala 50:65:@1306.4]
  assign _T_1958 = _T_1950[7]; // @[Bitwise.scala 50:65:@1307.4]
  assign _T_1959 = _T_1950[8]; // @[Bitwise.scala 50:65:@1308.4]
  assign _T_1960 = _T_1950[9]; // @[Bitwise.scala 50:65:@1309.4]
  assign _T_1961 = _T_1950[10]; // @[Bitwise.scala 50:65:@1310.4]
  assign _T_1962 = _T_1950[11]; // @[Bitwise.scala 50:65:@1311.4]
  assign _T_1963 = _T_1952 + _T_1953; // @[Bitwise.scala 48:55:@1312.4]
  assign _GEN_561 = {{1'd0}, _T_1951}; // @[Bitwise.scala 48:55:@1313.4]
  assign _T_1964 = _GEN_561 + _T_1963; // @[Bitwise.scala 48:55:@1313.4]
  assign _T_1965 = _T_1955 + _T_1956; // @[Bitwise.scala 48:55:@1314.4]
  assign _GEN_562 = {{1'd0}, _T_1954}; // @[Bitwise.scala 48:55:@1315.4]
  assign _T_1966 = _GEN_562 + _T_1965; // @[Bitwise.scala 48:55:@1315.4]
  assign _T_1967 = _T_1964 + _T_1966; // @[Bitwise.scala 48:55:@1316.4]
  assign _T_1968 = _T_1958 + _T_1959; // @[Bitwise.scala 48:55:@1317.4]
  assign _GEN_563 = {{1'd0}, _T_1957}; // @[Bitwise.scala 48:55:@1318.4]
  assign _T_1969 = _GEN_563 + _T_1968; // @[Bitwise.scala 48:55:@1318.4]
  assign _T_1970 = _T_1961 + _T_1962; // @[Bitwise.scala 48:55:@1319.4]
  assign _GEN_564 = {{1'd0}, _T_1960}; // @[Bitwise.scala 48:55:@1320.4]
  assign _T_1971 = _GEN_564 + _T_1970; // @[Bitwise.scala 48:55:@1320.4]
  assign _T_1972 = _T_1969 + _T_1971; // @[Bitwise.scala 48:55:@1321.4]
  assign _T_1973 = _T_1967 + _T_1972; // @[Bitwise.scala 48:55:@1322.4]
  assign _T_2037 = _T_1124[12:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1387.4]
  assign _T_2038 = _T_2037[0]; // @[Bitwise.scala 50:65:@1388.4]
  assign _T_2039 = _T_2037[1]; // @[Bitwise.scala 50:65:@1389.4]
  assign _T_2040 = _T_2037[2]; // @[Bitwise.scala 50:65:@1390.4]
  assign _T_2041 = _T_2037[3]; // @[Bitwise.scala 50:65:@1391.4]
  assign _T_2042 = _T_2037[4]; // @[Bitwise.scala 50:65:@1392.4]
  assign _T_2043 = _T_2037[5]; // @[Bitwise.scala 50:65:@1393.4]
  assign _T_2044 = _T_2037[6]; // @[Bitwise.scala 50:65:@1394.4]
  assign _T_2045 = _T_2037[7]; // @[Bitwise.scala 50:65:@1395.4]
  assign _T_2046 = _T_2037[8]; // @[Bitwise.scala 50:65:@1396.4]
  assign _T_2047 = _T_2037[9]; // @[Bitwise.scala 50:65:@1397.4]
  assign _T_2048 = _T_2037[10]; // @[Bitwise.scala 50:65:@1398.4]
  assign _T_2049 = _T_2037[11]; // @[Bitwise.scala 50:65:@1399.4]
  assign _T_2050 = _T_2037[12]; // @[Bitwise.scala 50:65:@1400.4]
  assign _T_2051 = _T_2039 + _T_2040; // @[Bitwise.scala 48:55:@1401.4]
  assign _GEN_565 = {{1'd0}, _T_2038}; // @[Bitwise.scala 48:55:@1402.4]
  assign _T_2052 = _GEN_565 + _T_2051; // @[Bitwise.scala 48:55:@1402.4]
  assign _T_2053 = _T_2042 + _T_2043; // @[Bitwise.scala 48:55:@1403.4]
  assign _GEN_566 = {{1'd0}, _T_2041}; // @[Bitwise.scala 48:55:@1404.4]
  assign _T_2054 = _GEN_566 + _T_2053; // @[Bitwise.scala 48:55:@1404.4]
  assign _T_2055 = _T_2052 + _T_2054; // @[Bitwise.scala 48:55:@1405.4]
  assign _T_2056 = _T_2045 + _T_2046; // @[Bitwise.scala 48:55:@1406.4]
  assign _GEN_567 = {{1'd0}, _T_2044}; // @[Bitwise.scala 48:55:@1407.4]
  assign _T_2057 = _GEN_567 + _T_2056; // @[Bitwise.scala 48:55:@1407.4]
  assign _T_2058 = _T_2047 + _T_2048; // @[Bitwise.scala 48:55:@1408.4]
  assign _T_2059 = _T_2049 + _T_2050; // @[Bitwise.scala 48:55:@1409.4]
  assign _T_2060 = _T_2058 + _T_2059; // @[Bitwise.scala 48:55:@1410.4]
  assign _T_2061 = _T_2057 + _T_2060; // @[Bitwise.scala 48:55:@1411.4]
  assign _T_2062 = _T_2055 + _T_2061; // @[Bitwise.scala 48:55:@1412.4]
  assign _T_2126 = _T_1124[13:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1477.4]
  assign _T_2127 = _T_2126[0]; // @[Bitwise.scala 50:65:@1478.4]
  assign _T_2128 = _T_2126[1]; // @[Bitwise.scala 50:65:@1479.4]
  assign _T_2129 = _T_2126[2]; // @[Bitwise.scala 50:65:@1480.4]
  assign _T_2130 = _T_2126[3]; // @[Bitwise.scala 50:65:@1481.4]
  assign _T_2131 = _T_2126[4]; // @[Bitwise.scala 50:65:@1482.4]
  assign _T_2132 = _T_2126[5]; // @[Bitwise.scala 50:65:@1483.4]
  assign _T_2133 = _T_2126[6]; // @[Bitwise.scala 50:65:@1484.4]
  assign _T_2134 = _T_2126[7]; // @[Bitwise.scala 50:65:@1485.4]
  assign _T_2135 = _T_2126[8]; // @[Bitwise.scala 50:65:@1486.4]
  assign _T_2136 = _T_2126[9]; // @[Bitwise.scala 50:65:@1487.4]
  assign _T_2137 = _T_2126[10]; // @[Bitwise.scala 50:65:@1488.4]
  assign _T_2138 = _T_2126[11]; // @[Bitwise.scala 50:65:@1489.4]
  assign _T_2139 = _T_2126[12]; // @[Bitwise.scala 50:65:@1490.4]
  assign _T_2140 = _T_2126[13]; // @[Bitwise.scala 50:65:@1491.4]
  assign _T_2141 = _T_2128 + _T_2129; // @[Bitwise.scala 48:55:@1492.4]
  assign _GEN_568 = {{1'd0}, _T_2127}; // @[Bitwise.scala 48:55:@1493.4]
  assign _T_2142 = _GEN_568 + _T_2141; // @[Bitwise.scala 48:55:@1493.4]
  assign _T_2143 = _T_2130 + _T_2131; // @[Bitwise.scala 48:55:@1494.4]
  assign _T_2144 = _T_2132 + _T_2133; // @[Bitwise.scala 48:55:@1495.4]
  assign _T_2145 = _T_2143 + _T_2144; // @[Bitwise.scala 48:55:@1496.4]
  assign _T_2146 = _T_2142 + _T_2145; // @[Bitwise.scala 48:55:@1497.4]
  assign _T_2147 = _T_2135 + _T_2136; // @[Bitwise.scala 48:55:@1498.4]
  assign _GEN_569 = {{1'd0}, _T_2134}; // @[Bitwise.scala 48:55:@1499.4]
  assign _T_2148 = _GEN_569 + _T_2147; // @[Bitwise.scala 48:55:@1499.4]
  assign _T_2149 = _T_2137 + _T_2138; // @[Bitwise.scala 48:55:@1500.4]
  assign _T_2150 = _T_2139 + _T_2140; // @[Bitwise.scala 48:55:@1501.4]
  assign _T_2151 = _T_2149 + _T_2150; // @[Bitwise.scala 48:55:@1502.4]
  assign _T_2152 = _T_2148 + _T_2151; // @[Bitwise.scala 48:55:@1503.4]
  assign _T_2153 = _T_2146 + _T_2152; // @[Bitwise.scala 48:55:@1504.4]
  assign _T_2217 = _T_1124[14:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1569.4]
  assign _T_2218 = _T_2217[0]; // @[Bitwise.scala 50:65:@1570.4]
  assign _T_2219 = _T_2217[1]; // @[Bitwise.scala 50:65:@1571.4]
  assign _T_2220 = _T_2217[2]; // @[Bitwise.scala 50:65:@1572.4]
  assign _T_2221 = _T_2217[3]; // @[Bitwise.scala 50:65:@1573.4]
  assign _T_2222 = _T_2217[4]; // @[Bitwise.scala 50:65:@1574.4]
  assign _T_2223 = _T_2217[5]; // @[Bitwise.scala 50:65:@1575.4]
  assign _T_2224 = _T_2217[6]; // @[Bitwise.scala 50:65:@1576.4]
  assign _T_2225 = _T_2217[7]; // @[Bitwise.scala 50:65:@1577.4]
  assign _T_2226 = _T_2217[8]; // @[Bitwise.scala 50:65:@1578.4]
  assign _T_2227 = _T_2217[9]; // @[Bitwise.scala 50:65:@1579.4]
  assign _T_2228 = _T_2217[10]; // @[Bitwise.scala 50:65:@1580.4]
  assign _T_2229 = _T_2217[11]; // @[Bitwise.scala 50:65:@1581.4]
  assign _T_2230 = _T_2217[12]; // @[Bitwise.scala 50:65:@1582.4]
  assign _T_2231 = _T_2217[13]; // @[Bitwise.scala 50:65:@1583.4]
  assign _T_2232 = _T_2217[14]; // @[Bitwise.scala 50:65:@1584.4]
  assign _T_2233 = _T_2219 + _T_2220; // @[Bitwise.scala 48:55:@1585.4]
  assign _GEN_570 = {{1'd0}, _T_2218}; // @[Bitwise.scala 48:55:@1586.4]
  assign _T_2234 = _GEN_570 + _T_2233; // @[Bitwise.scala 48:55:@1586.4]
  assign _T_2235 = _T_2221 + _T_2222; // @[Bitwise.scala 48:55:@1587.4]
  assign _T_2236 = _T_2223 + _T_2224; // @[Bitwise.scala 48:55:@1588.4]
  assign _T_2237 = _T_2235 + _T_2236; // @[Bitwise.scala 48:55:@1589.4]
  assign _T_2238 = _T_2234 + _T_2237; // @[Bitwise.scala 48:55:@1590.4]
  assign _T_2239 = _T_2225 + _T_2226; // @[Bitwise.scala 48:55:@1591.4]
  assign _T_2240 = _T_2227 + _T_2228; // @[Bitwise.scala 48:55:@1592.4]
  assign _T_2241 = _T_2239 + _T_2240; // @[Bitwise.scala 48:55:@1593.4]
  assign _T_2242 = _T_2229 + _T_2230; // @[Bitwise.scala 48:55:@1594.4]
  assign _T_2243 = _T_2231 + _T_2232; // @[Bitwise.scala 48:55:@1595.4]
  assign _T_2244 = _T_2242 + _T_2243; // @[Bitwise.scala 48:55:@1596.4]
  assign _T_2245 = _T_2241 + _T_2244; // @[Bitwise.scala 48:55:@1597.4]
  assign _T_2246 = _T_2238 + _T_2245; // @[Bitwise.scala 48:55:@1598.4]
  assign _T_2310 = _T_1124[15:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1663.4]
  assign _T_2311 = _T_2310[0]; // @[Bitwise.scala 50:65:@1664.4]
  assign _T_2312 = _T_2310[1]; // @[Bitwise.scala 50:65:@1665.4]
  assign _T_2313 = _T_2310[2]; // @[Bitwise.scala 50:65:@1666.4]
  assign _T_2314 = _T_2310[3]; // @[Bitwise.scala 50:65:@1667.4]
  assign _T_2315 = _T_2310[4]; // @[Bitwise.scala 50:65:@1668.4]
  assign _T_2316 = _T_2310[5]; // @[Bitwise.scala 50:65:@1669.4]
  assign _T_2317 = _T_2310[6]; // @[Bitwise.scala 50:65:@1670.4]
  assign _T_2318 = _T_2310[7]; // @[Bitwise.scala 50:65:@1671.4]
  assign _T_2319 = _T_2310[8]; // @[Bitwise.scala 50:65:@1672.4]
  assign _T_2320 = _T_2310[9]; // @[Bitwise.scala 50:65:@1673.4]
  assign _T_2321 = _T_2310[10]; // @[Bitwise.scala 50:65:@1674.4]
  assign _T_2322 = _T_2310[11]; // @[Bitwise.scala 50:65:@1675.4]
  assign _T_2323 = _T_2310[12]; // @[Bitwise.scala 50:65:@1676.4]
  assign _T_2324 = _T_2310[13]; // @[Bitwise.scala 50:65:@1677.4]
  assign _T_2325 = _T_2310[14]; // @[Bitwise.scala 50:65:@1678.4]
  assign _T_2326 = _T_2310[15]; // @[Bitwise.scala 50:65:@1679.4]
  assign _T_2327 = _T_2311 + _T_2312; // @[Bitwise.scala 48:55:@1680.4]
  assign _T_2328 = _T_2313 + _T_2314; // @[Bitwise.scala 48:55:@1681.4]
  assign _T_2329 = _T_2327 + _T_2328; // @[Bitwise.scala 48:55:@1682.4]
  assign _T_2330 = _T_2315 + _T_2316; // @[Bitwise.scala 48:55:@1683.4]
  assign _T_2331 = _T_2317 + _T_2318; // @[Bitwise.scala 48:55:@1684.4]
  assign _T_2332 = _T_2330 + _T_2331; // @[Bitwise.scala 48:55:@1685.4]
  assign _T_2333 = _T_2329 + _T_2332; // @[Bitwise.scala 48:55:@1686.4]
  assign _T_2334 = _T_2319 + _T_2320; // @[Bitwise.scala 48:55:@1687.4]
  assign _T_2335 = _T_2321 + _T_2322; // @[Bitwise.scala 48:55:@1688.4]
  assign _T_2336 = _T_2334 + _T_2335; // @[Bitwise.scala 48:55:@1689.4]
  assign _T_2337 = _T_2323 + _T_2324; // @[Bitwise.scala 48:55:@1690.4]
  assign _T_2338 = _T_2325 + _T_2326; // @[Bitwise.scala 48:55:@1691.4]
  assign _T_2339 = _T_2337 + _T_2338; // @[Bitwise.scala 48:55:@1692.4]
  assign _T_2340 = _T_2336 + _T_2339; // @[Bitwise.scala 48:55:@1693.4]
  assign _T_2341 = _T_2333 + _T_2340; // @[Bitwise.scala 48:55:@1694.4]
  assign _T_2405 = _T_1124[16:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1759.4]
  assign _T_2406 = _T_2405[0]; // @[Bitwise.scala 50:65:@1760.4]
  assign _T_2407 = _T_2405[1]; // @[Bitwise.scala 50:65:@1761.4]
  assign _T_2408 = _T_2405[2]; // @[Bitwise.scala 50:65:@1762.4]
  assign _T_2409 = _T_2405[3]; // @[Bitwise.scala 50:65:@1763.4]
  assign _T_2410 = _T_2405[4]; // @[Bitwise.scala 50:65:@1764.4]
  assign _T_2411 = _T_2405[5]; // @[Bitwise.scala 50:65:@1765.4]
  assign _T_2412 = _T_2405[6]; // @[Bitwise.scala 50:65:@1766.4]
  assign _T_2413 = _T_2405[7]; // @[Bitwise.scala 50:65:@1767.4]
  assign _T_2414 = _T_2405[8]; // @[Bitwise.scala 50:65:@1768.4]
  assign _T_2415 = _T_2405[9]; // @[Bitwise.scala 50:65:@1769.4]
  assign _T_2416 = _T_2405[10]; // @[Bitwise.scala 50:65:@1770.4]
  assign _T_2417 = _T_2405[11]; // @[Bitwise.scala 50:65:@1771.4]
  assign _T_2418 = _T_2405[12]; // @[Bitwise.scala 50:65:@1772.4]
  assign _T_2419 = _T_2405[13]; // @[Bitwise.scala 50:65:@1773.4]
  assign _T_2420 = _T_2405[14]; // @[Bitwise.scala 50:65:@1774.4]
  assign _T_2421 = _T_2405[15]; // @[Bitwise.scala 50:65:@1775.4]
  assign _T_2422 = _T_2405[16]; // @[Bitwise.scala 50:65:@1776.4]
  assign _T_2423 = _T_2406 + _T_2407; // @[Bitwise.scala 48:55:@1777.4]
  assign _T_2424 = _T_2408 + _T_2409; // @[Bitwise.scala 48:55:@1778.4]
  assign _T_2425 = _T_2423 + _T_2424; // @[Bitwise.scala 48:55:@1779.4]
  assign _T_2426 = _T_2410 + _T_2411; // @[Bitwise.scala 48:55:@1780.4]
  assign _T_2427 = _T_2412 + _T_2413; // @[Bitwise.scala 48:55:@1781.4]
  assign _T_2428 = _T_2426 + _T_2427; // @[Bitwise.scala 48:55:@1782.4]
  assign _T_2429 = _T_2425 + _T_2428; // @[Bitwise.scala 48:55:@1783.4]
  assign _T_2430 = _T_2414 + _T_2415; // @[Bitwise.scala 48:55:@1784.4]
  assign _T_2431 = _T_2416 + _T_2417; // @[Bitwise.scala 48:55:@1785.4]
  assign _T_2432 = _T_2430 + _T_2431; // @[Bitwise.scala 48:55:@1786.4]
  assign _T_2433 = _T_2418 + _T_2419; // @[Bitwise.scala 48:55:@1787.4]
  assign _T_2434 = _T_2421 + _T_2422; // @[Bitwise.scala 48:55:@1788.4]
  assign _GEN_571 = {{1'd0}, _T_2420}; // @[Bitwise.scala 48:55:@1789.4]
  assign _T_2435 = _GEN_571 + _T_2434; // @[Bitwise.scala 48:55:@1789.4]
  assign _GEN_572 = {{1'd0}, _T_2433}; // @[Bitwise.scala 48:55:@1790.4]
  assign _T_2436 = _GEN_572 + _T_2435; // @[Bitwise.scala 48:55:@1790.4]
  assign _GEN_573 = {{1'd0}, _T_2432}; // @[Bitwise.scala 48:55:@1791.4]
  assign _T_2437 = _GEN_573 + _T_2436; // @[Bitwise.scala 48:55:@1791.4]
  assign _GEN_574 = {{1'd0}, _T_2429}; // @[Bitwise.scala 48:55:@1792.4]
  assign _T_2438 = _GEN_574 + _T_2437; // @[Bitwise.scala 48:55:@1792.4]
  assign _T_2502 = _T_1124[17:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1857.4]
  assign _T_2503 = _T_2502[0]; // @[Bitwise.scala 50:65:@1858.4]
  assign _T_2504 = _T_2502[1]; // @[Bitwise.scala 50:65:@1859.4]
  assign _T_2505 = _T_2502[2]; // @[Bitwise.scala 50:65:@1860.4]
  assign _T_2506 = _T_2502[3]; // @[Bitwise.scala 50:65:@1861.4]
  assign _T_2507 = _T_2502[4]; // @[Bitwise.scala 50:65:@1862.4]
  assign _T_2508 = _T_2502[5]; // @[Bitwise.scala 50:65:@1863.4]
  assign _T_2509 = _T_2502[6]; // @[Bitwise.scala 50:65:@1864.4]
  assign _T_2510 = _T_2502[7]; // @[Bitwise.scala 50:65:@1865.4]
  assign _T_2511 = _T_2502[8]; // @[Bitwise.scala 50:65:@1866.4]
  assign _T_2512 = _T_2502[9]; // @[Bitwise.scala 50:65:@1867.4]
  assign _T_2513 = _T_2502[10]; // @[Bitwise.scala 50:65:@1868.4]
  assign _T_2514 = _T_2502[11]; // @[Bitwise.scala 50:65:@1869.4]
  assign _T_2515 = _T_2502[12]; // @[Bitwise.scala 50:65:@1870.4]
  assign _T_2516 = _T_2502[13]; // @[Bitwise.scala 50:65:@1871.4]
  assign _T_2517 = _T_2502[14]; // @[Bitwise.scala 50:65:@1872.4]
  assign _T_2518 = _T_2502[15]; // @[Bitwise.scala 50:65:@1873.4]
  assign _T_2519 = _T_2502[16]; // @[Bitwise.scala 50:65:@1874.4]
  assign _T_2520 = _T_2502[17]; // @[Bitwise.scala 50:65:@1875.4]
  assign _T_2521 = _T_2503 + _T_2504; // @[Bitwise.scala 48:55:@1876.4]
  assign _T_2522 = _T_2505 + _T_2506; // @[Bitwise.scala 48:55:@1877.4]
  assign _T_2523 = _T_2521 + _T_2522; // @[Bitwise.scala 48:55:@1878.4]
  assign _T_2524 = _T_2507 + _T_2508; // @[Bitwise.scala 48:55:@1879.4]
  assign _T_2525 = _T_2510 + _T_2511; // @[Bitwise.scala 48:55:@1880.4]
  assign _GEN_575 = {{1'd0}, _T_2509}; // @[Bitwise.scala 48:55:@1881.4]
  assign _T_2526 = _GEN_575 + _T_2525; // @[Bitwise.scala 48:55:@1881.4]
  assign _GEN_576 = {{1'd0}, _T_2524}; // @[Bitwise.scala 48:55:@1882.4]
  assign _T_2527 = _GEN_576 + _T_2526; // @[Bitwise.scala 48:55:@1882.4]
  assign _GEN_577 = {{1'd0}, _T_2523}; // @[Bitwise.scala 48:55:@1883.4]
  assign _T_2528 = _GEN_577 + _T_2527; // @[Bitwise.scala 48:55:@1883.4]
  assign _T_2529 = _T_2512 + _T_2513; // @[Bitwise.scala 48:55:@1884.4]
  assign _T_2530 = _T_2514 + _T_2515; // @[Bitwise.scala 48:55:@1885.4]
  assign _T_2531 = _T_2529 + _T_2530; // @[Bitwise.scala 48:55:@1886.4]
  assign _T_2532 = _T_2516 + _T_2517; // @[Bitwise.scala 48:55:@1887.4]
  assign _T_2533 = _T_2519 + _T_2520; // @[Bitwise.scala 48:55:@1888.4]
  assign _GEN_578 = {{1'd0}, _T_2518}; // @[Bitwise.scala 48:55:@1889.4]
  assign _T_2534 = _GEN_578 + _T_2533; // @[Bitwise.scala 48:55:@1889.4]
  assign _GEN_579 = {{1'd0}, _T_2532}; // @[Bitwise.scala 48:55:@1890.4]
  assign _T_2535 = _GEN_579 + _T_2534; // @[Bitwise.scala 48:55:@1890.4]
  assign _GEN_580 = {{1'd0}, _T_2531}; // @[Bitwise.scala 48:55:@1891.4]
  assign _T_2536 = _GEN_580 + _T_2535; // @[Bitwise.scala 48:55:@1891.4]
  assign _T_2537 = _T_2528 + _T_2536; // @[Bitwise.scala 48:55:@1892.4]
  assign _T_2601 = _T_1124[18:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@1957.4]
  assign _T_2602 = _T_2601[0]; // @[Bitwise.scala 50:65:@1958.4]
  assign _T_2603 = _T_2601[1]; // @[Bitwise.scala 50:65:@1959.4]
  assign _T_2604 = _T_2601[2]; // @[Bitwise.scala 50:65:@1960.4]
  assign _T_2605 = _T_2601[3]; // @[Bitwise.scala 50:65:@1961.4]
  assign _T_2606 = _T_2601[4]; // @[Bitwise.scala 50:65:@1962.4]
  assign _T_2607 = _T_2601[5]; // @[Bitwise.scala 50:65:@1963.4]
  assign _T_2608 = _T_2601[6]; // @[Bitwise.scala 50:65:@1964.4]
  assign _T_2609 = _T_2601[7]; // @[Bitwise.scala 50:65:@1965.4]
  assign _T_2610 = _T_2601[8]; // @[Bitwise.scala 50:65:@1966.4]
  assign _T_2611 = _T_2601[9]; // @[Bitwise.scala 50:65:@1967.4]
  assign _T_2612 = _T_2601[10]; // @[Bitwise.scala 50:65:@1968.4]
  assign _T_2613 = _T_2601[11]; // @[Bitwise.scala 50:65:@1969.4]
  assign _T_2614 = _T_2601[12]; // @[Bitwise.scala 50:65:@1970.4]
  assign _T_2615 = _T_2601[13]; // @[Bitwise.scala 50:65:@1971.4]
  assign _T_2616 = _T_2601[14]; // @[Bitwise.scala 50:65:@1972.4]
  assign _T_2617 = _T_2601[15]; // @[Bitwise.scala 50:65:@1973.4]
  assign _T_2618 = _T_2601[16]; // @[Bitwise.scala 50:65:@1974.4]
  assign _T_2619 = _T_2601[17]; // @[Bitwise.scala 50:65:@1975.4]
  assign _T_2620 = _T_2601[18]; // @[Bitwise.scala 50:65:@1976.4]
  assign _T_2621 = _T_2602 + _T_2603; // @[Bitwise.scala 48:55:@1977.4]
  assign _T_2622 = _T_2604 + _T_2605; // @[Bitwise.scala 48:55:@1978.4]
  assign _T_2623 = _T_2621 + _T_2622; // @[Bitwise.scala 48:55:@1979.4]
  assign _T_2624 = _T_2606 + _T_2607; // @[Bitwise.scala 48:55:@1980.4]
  assign _T_2625 = _T_2609 + _T_2610; // @[Bitwise.scala 48:55:@1981.4]
  assign _GEN_581 = {{1'd0}, _T_2608}; // @[Bitwise.scala 48:55:@1982.4]
  assign _T_2626 = _GEN_581 + _T_2625; // @[Bitwise.scala 48:55:@1982.4]
  assign _GEN_582 = {{1'd0}, _T_2624}; // @[Bitwise.scala 48:55:@1983.4]
  assign _T_2627 = _GEN_582 + _T_2626; // @[Bitwise.scala 48:55:@1983.4]
  assign _GEN_583 = {{1'd0}, _T_2623}; // @[Bitwise.scala 48:55:@1984.4]
  assign _T_2628 = _GEN_583 + _T_2627; // @[Bitwise.scala 48:55:@1984.4]
  assign _T_2629 = _T_2611 + _T_2612; // @[Bitwise.scala 48:55:@1985.4]
  assign _T_2630 = _T_2614 + _T_2615; // @[Bitwise.scala 48:55:@1986.4]
  assign _GEN_584 = {{1'd0}, _T_2613}; // @[Bitwise.scala 48:55:@1987.4]
  assign _T_2631 = _GEN_584 + _T_2630; // @[Bitwise.scala 48:55:@1987.4]
  assign _GEN_585 = {{1'd0}, _T_2629}; // @[Bitwise.scala 48:55:@1988.4]
  assign _T_2632 = _GEN_585 + _T_2631; // @[Bitwise.scala 48:55:@1988.4]
  assign _T_2633 = _T_2616 + _T_2617; // @[Bitwise.scala 48:55:@1989.4]
  assign _T_2634 = _T_2619 + _T_2620; // @[Bitwise.scala 48:55:@1990.4]
  assign _GEN_586 = {{1'd0}, _T_2618}; // @[Bitwise.scala 48:55:@1991.4]
  assign _T_2635 = _GEN_586 + _T_2634; // @[Bitwise.scala 48:55:@1991.4]
  assign _GEN_587 = {{1'd0}, _T_2633}; // @[Bitwise.scala 48:55:@1992.4]
  assign _T_2636 = _GEN_587 + _T_2635; // @[Bitwise.scala 48:55:@1992.4]
  assign _T_2637 = _T_2632 + _T_2636; // @[Bitwise.scala 48:55:@1993.4]
  assign _T_2638 = _T_2628 + _T_2637; // @[Bitwise.scala 48:55:@1994.4]
  assign _T_2702 = _T_1124[19:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2059.4]
  assign _T_2703 = _T_2702[0]; // @[Bitwise.scala 50:65:@2060.4]
  assign _T_2704 = _T_2702[1]; // @[Bitwise.scala 50:65:@2061.4]
  assign _T_2705 = _T_2702[2]; // @[Bitwise.scala 50:65:@2062.4]
  assign _T_2706 = _T_2702[3]; // @[Bitwise.scala 50:65:@2063.4]
  assign _T_2707 = _T_2702[4]; // @[Bitwise.scala 50:65:@2064.4]
  assign _T_2708 = _T_2702[5]; // @[Bitwise.scala 50:65:@2065.4]
  assign _T_2709 = _T_2702[6]; // @[Bitwise.scala 50:65:@2066.4]
  assign _T_2710 = _T_2702[7]; // @[Bitwise.scala 50:65:@2067.4]
  assign _T_2711 = _T_2702[8]; // @[Bitwise.scala 50:65:@2068.4]
  assign _T_2712 = _T_2702[9]; // @[Bitwise.scala 50:65:@2069.4]
  assign _T_2713 = _T_2702[10]; // @[Bitwise.scala 50:65:@2070.4]
  assign _T_2714 = _T_2702[11]; // @[Bitwise.scala 50:65:@2071.4]
  assign _T_2715 = _T_2702[12]; // @[Bitwise.scala 50:65:@2072.4]
  assign _T_2716 = _T_2702[13]; // @[Bitwise.scala 50:65:@2073.4]
  assign _T_2717 = _T_2702[14]; // @[Bitwise.scala 50:65:@2074.4]
  assign _T_2718 = _T_2702[15]; // @[Bitwise.scala 50:65:@2075.4]
  assign _T_2719 = _T_2702[16]; // @[Bitwise.scala 50:65:@2076.4]
  assign _T_2720 = _T_2702[17]; // @[Bitwise.scala 50:65:@2077.4]
  assign _T_2721 = _T_2702[18]; // @[Bitwise.scala 50:65:@2078.4]
  assign _T_2722 = _T_2702[19]; // @[Bitwise.scala 50:65:@2079.4]
  assign _T_2723 = _T_2703 + _T_2704; // @[Bitwise.scala 48:55:@2080.4]
  assign _T_2724 = _T_2706 + _T_2707; // @[Bitwise.scala 48:55:@2081.4]
  assign _GEN_588 = {{1'd0}, _T_2705}; // @[Bitwise.scala 48:55:@2082.4]
  assign _T_2725 = _GEN_588 + _T_2724; // @[Bitwise.scala 48:55:@2082.4]
  assign _GEN_589 = {{1'd0}, _T_2723}; // @[Bitwise.scala 48:55:@2083.4]
  assign _T_2726 = _GEN_589 + _T_2725; // @[Bitwise.scala 48:55:@2083.4]
  assign _T_2727 = _T_2708 + _T_2709; // @[Bitwise.scala 48:55:@2084.4]
  assign _T_2728 = _T_2711 + _T_2712; // @[Bitwise.scala 48:55:@2085.4]
  assign _GEN_590 = {{1'd0}, _T_2710}; // @[Bitwise.scala 48:55:@2086.4]
  assign _T_2729 = _GEN_590 + _T_2728; // @[Bitwise.scala 48:55:@2086.4]
  assign _GEN_591 = {{1'd0}, _T_2727}; // @[Bitwise.scala 48:55:@2087.4]
  assign _T_2730 = _GEN_591 + _T_2729; // @[Bitwise.scala 48:55:@2087.4]
  assign _T_2731 = _T_2726 + _T_2730; // @[Bitwise.scala 48:55:@2088.4]
  assign _T_2732 = _T_2713 + _T_2714; // @[Bitwise.scala 48:55:@2089.4]
  assign _T_2733 = _T_2716 + _T_2717; // @[Bitwise.scala 48:55:@2090.4]
  assign _GEN_592 = {{1'd0}, _T_2715}; // @[Bitwise.scala 48:55:@2091.4]
  assign _T_2734 = _GEN_592 + _T_2733; // @[Bitwise.scala 48:55:@2091.4]
  assign _GEN_593 = {{1'd0}, _T_2732}; // @[Bitwise.scala 48:55:@2092.4]
  assign _T_2735 = _GEN_593 + _T_2734; // @[Bitwise.scala 48:55:@2092.4]
  assign _T_2736 = _T_2718 + _T_2719; // @[Bitwise.scala 48:55:@2093.4]
  assign _T_2737 = _T_2721 + _T_2722; // @[Bitwise.scala 48:55:@2094.4]
  assign _GEN_594 = {{1'd0}, _T_2720}; // @[Bitwise.scala 48:55:@2095.4]
  assign _T_2738 = _GEN_594 + _T_2737; // @[Bitwise.scala 48:55:@2095.4]
  assign _GEN_595 = {{1'd0}, _T_2736}; // @[Bitwise.scala 48:55:@2096.4]
  assign _T_2739 = _GEN_595 + _T_2738; // @[Bitwise.scala 48:55:@2096.4]
  assign _T_2740 = _T_2735 + _T_2739; // @[Bitwise.scala 48:55:@2097.4]
  assign _T_2741 = _T_2731 + _T_2740; // @[Bitwise.scala 48:55:@2098.4]
  assign _T_2805 = _T_1124[20:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2163.4]
  assign _T_2806 = _T_2805[0]; // @[Bitwise.scala 50:65:@2164.4]
  assign _T_2807 = _T_2805[1]; // @[Bitwise.scala 50:65:@2165.4]
  assign _T_2808 = _T_2805[2]; // @[Bitwise.scala 50:65:@2166.4]
  assign _T_2809 = _T_2805[3]; // @[Bitwise.scala 50:65:@2167.4]
  assign _T_2810 = _T_2805[4]; // @[Bitwise.scala 50:65:@2168.4]
  assign _T_2811 = _T_2805[5]; // @[Bitwise.scala 50:65:@2169.4]
  assign _T_2812 = _T_2805[6]; // @[Bitwise.scala 50:65:@2170.4]
  assign _T_2813 = _T_2805[7]; // @[Bitwise.scala 50:65:@2171.4]
  assign _T_2814 = _T_2805[8]; // @[Bitwise.scala 50:65:@2172.4]
  assign _T_2815 = _T_2805[9]; // @[Bitwise.scala 50:65:@2173.4]
  assign _T_2816 = _T_2805[10]; // @[Bitwise.scala 50:65:@2174.4]
  assign _T_2817 = _T_2805[11]; // @[Bitwise.scala 50:65:@2175.4]
  assign _T_2818 = _T_2805[12]; // @[Bitwise.scala 50:65:@2176.4]
  assign _T_2819 = _T_2805[13]; // @[Bitwise.scala 50:65:@2177.4]
  assign _T_2820 = _T_2805[14]; // @[Bitwise.scala 50:65:@2178.4]
  assign _T_2821 = _T_2805[15]; // @[Bitwise.scala 50:65:@2179.4]
  assign _T_2822 = _T_2805[16]; // @[Bitwise.scala 50:65:@2180.4]
  assign _T_2823 = _T_2805[17]; // @[Bitwise.scala 50:65:@2181.4]
  assign _T_2824 = _T_2805[18]; // @[Bitwise.scala 50:65:@2182.4]
  assign _T_2825 = _T_2805[19]; // @[Bitwise.scala 50:65:@2183.4]
  assign _T_2826 = _T_2805[20]; // @[Bitwise.scala 50:65:@2184.4]
  assign _T_2827 = _T_2806 + _T_2807; // @[Bitwise.scala 48:55:@2185.4]
  assign _T_2828 = _T_2809 + _T_2810; // @[Bitwise.scala 48:55:@2186.4]
  assign _GEN_596 = {{1'd0}, _T_2808}; // @[Bitwise.scala 48:55:@2187.4]
  assign _T_2829 = _GEN_596 + _T_2828; // @[Bitwise.scala 48:55:@2187.4]
  assign _GEN_597 = {{1'd0}, _T_2827}; // @[Bitwise.scala 48:55:@2188.4]
  assign _T_2830 = _GEN_597 + _T_2829; // @[Bitwise.scala 48:55:@2188.4]
  assign _T_2831 = _T_2811 + _T_2812; // @[Bitwise.scala 48:55:@2189.4]
  assign _T_2832 = _T_2814 + _T_2815; // @[Bitwise.scala 48:55:@2190.4]
  assign _GEN_598 = {{1'd0}, _T_2813}; // @[Bitwise.scala 48:55:@2191.4]
  assign _T_2833 = _GEN_598 + _T_2832; // @[Bitwise.scala 48:55:@2191.4]
  assign _GEN_599 = {{1'd0}, _T_2831}; // @[Bitwise.scala 48:55:@2192.4]
  assign _T_2834 = _GEN_599 + _T_2833; // @[Bitwise.scala 48:55:@2192.4]
  assign _T_2835 = _T_2830 + _T_2834; // @[Bitwise.scala 48:55:@2193.4]
  assign _T_2836 = _T_2816 + _T_2817; // @[Bitwise.scala 48:55:@2194.4]
  assign _T_2837 = _T_2819 + _T_2820; // @[Bitwise.scala 48:55:@2195.4]
  assign _GEN_600 = {{1'd0}, _T_2818}; // @[Bitwise.scala 48:55:@2196.4]
  assign _T_2838 = _GEN_600 + _T_2837; // @[Bitwise.scala 48:55:@2196.4]
  assign _GEN_601 = {{1'd0}, _T_2836}; // @[Bitwise.scala 48:55:@2197.4]
  assign _T_2839 = _GEN_601 + _T_2838; // @[Bitwise.scala 48:55:@2197.4]
  assign _T_2840 = _T_2822 + _T_2823; // @[Bitwise.scala 48:55:@2198.4]
  assign _GEN_602 = {{1'd0}, _T_2821}; // @[Bitwise.scala 48:55:@2199.4]
  assign _T_2841 = _GEN_602 + _T_2840; // @[Bitwise.scala 48:55:@2199.4]
  assign _T_2842 = _T_2825 + _T_2826; // @[Bitwise.scala 48:55:@2200.4]
  assign _GEN_603 = {{1'd0}, _T_2824}; // @[Bitwise.scala 48:55:@2201.4]
  assign _T_2843 = _GEN_603 + _T_2842; // @[Bitwise.scala 48:55:@2201.4]
  assign _T_2844 = _T_2841 + _T_2843; // @[Bitwise.scala 48:55:@2202.4]
  assign _T_2845 = _T_2839 + _T_2844; // @[Bitwise.scala 48:55:@2203.4]
  assign _T_2846 = _T_2835 + _T_2845; // @[Bitwise.scala 48:55:@2204.4]
  assign _T_2910 = _T_1124[21:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2269.4]
  assign _T_2911 = _T_2910[0]; // @[Bitwise.scala 50:65:@2270.4]
  assign _T_2912 = _T_2910[1]; // @[Bitwise.scala 50:65:@2271.4]
  assign _T_2913 = _T_2910[2]; // @[Bitwise.scala 50:65:@2272.4]
  assign _T_2914 = _T_2910[3]; // @[Bitwise.scala 50:65:@2273.4]
  assign _T_2915 = _T_2910[4]; // @[Bitwise.scala 50:65:@2274.4]
  assign _T_2916 = _T_2910[5]; // @[Bitwise.scala 50:65:@2275.4]
  assign _T_2917 = _T_2910[6]; // @[Bitwise.scala 50:65:@2276.4]
  assign _T_2918 = _T_2910[7]; // @[Bitwise.scala 50:65:@2277.4]
  assign _T_2919 = _T_2910[8]; // @[Bitwise.scala 50:65:@2278.4]
  assign _T_2920 = _T_2910[9]; // @[Bitwise.scala 50:65:@2279.4]
  assign _T_2921 = _T_2910[10]; // @[Bitwise.scala 50:65:@2280.4]
  assign _T_2922 = _T_2910[11]; // @[Bitwise.scala 50:65:@2281.4]
  assign _T_2923 = _T_2910[12]; // @[Bitwise.scala 50:65:@2282.4]
  assign _T_2924 = _T_2910[13]; // @[Bitwise.scala 50:65:@2283.4]
  assign _T_2925 = _T_2910[14]; // @[Bitwise.scala 50:65:@2284.4]
  assign _T_2926 = _T_2910[15]; // @[Bitwise.scala 50:65:@2285.4]
  assign _T_2927 = _T_2910[16]; // @[Bitwise.scala 50:65:@2286.4]
  assign _T_2928 = _T_2910[17]; // @[Bitwise.scala 50:65:@2287.4]
  assign _T_2929 = _T_2910[18]; // @[Bitwise.scala 50:65:@2288.4]
  assign _T_2930 = _T_2910[19]; // @[Bitwise.scala 50:65:@2289.4]
  assign _T_2931 = _T_2910[20]; // @[Bitwise.scala 50:65:@2290.4]
  assign _T_2932 = _T_2910[21]; // @[Bitwise.scala 50:65:@2291.4]
  assign _T_2933 = _T_2911 + _T_2912; // @[Bitwise.scala 48:55:@2292.4]
  assign _T_2934 = _T_2914 + _T_2915; // @[Bitwise.scala 48:55:@2293.4]
  assign _GEN_604 = {{1'd0}, _T_2913}; // @[Bitwise.scala 48:55:@2294.4]
  assign _T_2935 = _GEN_604 + _T_2934; // @[Bitwise.scala 48:55:@2294.4]
  assign _GEN_605 = {{1'd0}, _T_2933}; // @[Bitwise.scala 48:55:@2295.4]
  assign _T_2936 = _GEN_605 + _T_2935; // @[Bitwise.scala 48:55:@2295.4]
  assign _T_2937 = _T_2917 + _T_2918; // @[Bitwise.scala 48:55:@2296.4]
  assign _GEN_606 = {{1'd0}, _T_2916}; // @[Bitwise.scala 48:55:@2297.4]
  assign _T_2938 = _GEN_606 + _T_2937; // @[Bitwise.scala 48:55:@2297.4]
  assign _T_2939 = _T_2920 + _T_2921; // @[Bitwise.scala 48:55:@2298.4]
  assign _GEN_607 = {{1'd0}, _T_2919}; // @[Bitwise.scala 48:55:@2299.4]
  assign _T_2940 = _GEN_607 + _T_2939; // @[Bitwise.scala 48:55:@2299.4]
  assign _T_2941 = _T_2938 + _T_2940; // @[Bitwise.scala 48:55:@2300.4]
  assign _T_2942 = _T_2936 + _T_2941; // @[Bitwise.scala 48:55:@2301.4]
  assign _T_2943 = _T_2922 + _T_2923; // @[Bitwise.scala 48:55:@2302.4]
  assign _T_2944 = _T_2925 + _T_2926; // @[Bitwise.scala 48:55:@2303.4]
  assign _GEN_608 = {{1'd0}, _T_2924}; // @[Bitwise.scala 48:55:@2304.4]
  assign _T_2945 = _GEN_608 + _T_2944; // @[Bitwise.scala 48:55:@2304.4]
  assign _GEN_609 = {{1'd0}, _T_2943}; // @[Bitwise.scala 48:55:@2305.4]
  assign _T_2946 = _GEN_609 + _T_2945; // @[Bitwise.scala 48:55:@2305.4]
  assign _T_2947 = _T_2928 + _T_2929; // @[Bitwise.scala 48:55:@2306.4]
  assign _GEN_610 = {{1'd0}, _T_2927}; // @[Bitwise.scala 48:55:@2307.4]
  assign _T_2948 = _GEN_610 + _T_2947; // @[Bitwise.scala 48:55:@2307.4]
  assign _T_2949 = _T_2931 + _T_2932; // @[Bitwise.scala 48:55:@2308.4]
  assign _GEN_611 = {{1'd0}, _T_2930}; // @[Bitwise.scala 48:55:@2309.4]
  assign _T_2950 = _GEN_611 + _T_2949; // @[Bitwise.scala 48:55:@2309.4]
  assign _T_2951 = _T_2948 + _T_2950; // @[Bitwise.scala 48:55:@2310.4]
  assign _T_2952 = _T_2946 + _T_2951; // @[Bitwise.scala 48:55:@2311.4]
  assign _T_2953 = _T_2942 + _T_2952; // @[Bitwise.scala 48:55:@2312.4]
  assign _T_3017 = _T_1124[22:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2377.4]
  assign _T_3018 = _T_3017[0]; // @[Bitwise.scala 50:65:@2378.4]
  assign _T_3019 = _T_3017[1]; // @[Bitwise.scala 50:65:@2379.4]
  assign _T_3020 = _T_3017[2]; // @[Bitwise.scala 50:65:@2380.4]
  assign _T_3021 = _T_3017[3]; // @[Bitwise.scala 50:65:@2381.4]
  assign _T_3022 = _T_3017[4]; // @[Bitwise.scala 50:65:@2382.4]
  assign _T_3023 = _T_3017[5]; // @[Bitwise.scala 50:65:@2383.4]
  assign _T_3024 = _T_3017[6]; // @[Bitwise.scala 50:65:@2384.4]
  assign _T_3025 = _T_3017[7]; // @[Bitwise.scala 50:65:@2385.4]
  assign _T_3026 = _T_3017[8]; // @[Bitwise.scala 50:65:@2386.4]
  assign _T_3027 = _T_3017[9]; // @[Bitwise.scala 50:65:@2387.4]
  assign _T_3028 = _T_3017[10]; // @[Bitwise.scala 50:65:@2388.4]
  assign _T_3029 = _T_3017[11]; // @[Bitwise.scala 50:65:@2389.4]
  assign _T_3030 = _T_3017[12]; // @[Bitwise.scala 50:65:@2390.4]
  assign _T_3031 = _T_3017[13]; // @[Bitwise.scala 50:65:@2391.4]
  assign _T_3032 = _T_3017[14]; // @[Bitwise.scala 50:65:@2392.4]
  assign _T_3033 = _T_3017[15]; // @[Bitwise.scala 50:65:@2393.4]
  assign _T_3034 = _T_3017[16]; // @[Bitwise.scala 50:65:@2394.4]
  assign _T_3035 = _T_3017[17]; // @[Bitwise.scala 50:65:@2395.4]
  assign _T_3036 = _T_3017[18]; // @[Bitwise.scala 50:65:@2396.4]
  assign _T_3037 = _T_3017[19]; // @[Bitwise.scala 50:65:@2397.4]
  assign _T_3038 = _T_3017[20]; // @[Bitwise.scala 50:65:@2398.4]
  assign _T_3039 = _T_3017[21]; // @[Bitwise.scala 50:65:@2399.4]
  assign _T_3040 = _T_3017[22]; // @[Bitwise.scala 50:65:@2400.4]
  assign _T_3041 = _T_3018 + _T_3019; // @[Bitwise.scala 48:55:@2401.4]
  assign _T_3042 = _T_3021 + _T_3022; // @[Bitwise.scala 48:55:@2402.4]
  assign _GEN_612 = {{1'd0}, _T_3020}; // @[Bitwise.scala 48:55:@2403.4]
  assign _T_3043 = _GEN_612 + _T_3042; // @[Bitwise.scala 48:55:@2403.4]
  assign _GEN_613 = {{1'd0}, _T_3041}; // @[Bitwise.scala 48:55:@2404.4]
  assign _T_3044 = _GEN_613 + _T_3043; // @[Bitwise.scala 48:55:@2404.4]
  assign _T_3045 = _T_3024 + _T_3025; // @[Bitwise.scala 48:55:@2405.4]
  assign _GEN_614 = {{1'd0}, _T_3023}; // @[Bitwise.scala 48:55:@2406.4]
  assign _T_3046 = _GEN_614 + _T_3045; // @[Bitwise.scala 48:55:@2406.4]
  assign _T_3047 = _T_3027 + _T_3028; // @[Bitwise.scala 48:55:@2407.4]
  assign _GEN_615 = {{1'd0}, _T_3026}; // @[Bitwise.scala 48:55:@2408.4]
  assign _T_3048 = _GEN_615 + _T_3047; // @[Bitwise.scala 48:55:@2408.4]
  assign _T_3049 = _T_3046 + _T_3048; // @[Bitwise.scala 48:55:@2409.4]
  assign _T_3050 = _T_3044 + _T_3049; // @[Bitwise.scala 48:55:@2410.4]
  assign _T_3051 = _T_3030 + _T_3031; // @[Bitwise.scala 48:55:@2411.4]
  assign _GEN_616 = {{1'd0}, _T_3029}; // @[Bitwise.scala 48:55:@2412.4]
  assign _T_3052 = _GEN_616 + _T_3051; // @[Bitwise.scala 48:55:@2412.4]
  assign _T_3053 = _T_3033 + _T_3034; // @[Bitwise.scala 48:55:@2413.4]
  assign _GEN_617 = {{1'd0}, _T_3032}; // @[Bitwise.scala 48:55:@2414.4]
  assign _T_3054 = _GEN_617 + _T_3053; // @[Bitwise.scala 48:55:@2414.4]
  assign _T_3055 = _T_3052 + _T_3054; // @[Bitwise.scala 48:55:@2415.4]
  assign _T_3056 = _T_3036 + _T_3037; // @[Bitwise.scala 48:55:@2416.4]
  assign _GEN_618 = {{1'd0}, _T_3035}; // @[Bitwise.scala 48:55:@2417.4]
  assign _T_3057 = _GEN_618 + _T_3056; // @[Bitwise.scala 48:55:@2417.4]
  assign _T_3058 = _T_3039 + _T_3040; // @[Bitwise.scala 48:55:@2418.4]
  assign _GEN_619 = {{1'd0}, _T_3038}; // @[Bitwise.scala 48:55:@2419.4]
  assign _T_3059 = _GEN_619 + _T_3058; // @[Bitwise.scala 48:55:@2419.4]
  assign _T_3060 = _T_3057 + _T_3059; // @[Bitwise.scala 48:55:@2420.4]
  assign _T_3061 = _T_3055 + _T_3060; // @[Bitwise.scala 48:55:@2421.4]
  assign _T_3062 = _T_3050 + _T_3061; // @[Bitwise.scala 48:55:@2422.4]
  assign _T_3126 = _T_1124[23:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2487.4]
  assign _T_3127 = _T_3126[0]; // @[Bitwise.scala 50:65:@2488.4]
  assign _T_3128 = _T_3126[1]; // @[Bitwise.scala 50:65:@2489.4]
  assign _T_3129 = _T_3126[2]; // @[Bitwise.scala 50:65:@2490.4]
  assign _T_3130 = _T_3126[3]; // @[Bitwise.scala 50:65:@2491.4]
  assign _T_3131 = _T_3126[4]; // @[Bitwise.scala 50:65:@2492.4]
  assign _T_3132 = _T_3126[5]; // @[Bitwise.scala 50:65:@2493.4]
  assign _T_3133 = _T_3126[6]; // @[Bitwise.scala 50:65:@2494.4]
  assign _T_3134 = _T_3126[7]; // @[Bitwise.scala 50:65:@2495.4]
  assign _T_3135 = _T_3126[8]; // @[Bitwise.scala 50:65:@2496.4]
  assign _T_3136 = _T_3126[9]; // @[Bitwise.scala 50:65:@2497.4]
  assign _T_3137 = _T_3126[10]; // @[Bitwise.scala 50:65:@2498.4]
  assign _T_3138 = _T_3126[11]; // @[Bitwise.scala 50:65:@2499.4]
  assign _T_3139 = _T_3126[12]; // @[Bitwise.scala 50:65:@2500.4]
  assign _T_3140 = _T_3126[13]; // @[Bitwise.scala 50:65:@2501.4]
  assign _T_3141 = _T_3126[14]; // @[Bitwise.scala 50:65:@2502.4]
  assign _T_3142 = _T_3126[15]; // @[Bitwise.scala 50:65:@2503.4]
  assign _T_3143 = _T_3126[16]; // @[Bitwise.scala 50:65:@2504.4]
  assign _T_3144 = _T_3126[17]; // @[Bitwise.scala 50:65:@2505.4]
  assign _T_3145 = _T_3126[18]; // @[Bitwise.scala 50:65:@2506.4]
  assign _T_3146 = _T_3126[19]; // @[Bitwise.scala 50:65:@2507.4]
  assign _T_3147 = _T_3126[20]; // @[Bitwise.scala 50:65:@2508.4]
  assign _T_3148 = _T_3126[21]; // @[Bitwise.scala 50:65:@2509.4]
  assign _T_3149 = _T_3126[22]; // @[Bitwise.scala 50:65:@2510.4]
  assign _T_3150 = _T_3126[23]; // @[Bitwise.scala 50:65:@2511.4]
  assign _T_3151 = _T_3128 + _T_3129; // @[Bitwise.scala 48:55:@2512.4]
  assign _GEN_620 = {{1'd0}, _T_3127}; // @[Bitwise.scala 48:55:@2513.4]
  assign _T_3152 = _GEN_620 + _T_3151; // @[Bitwise.scala 48:55:@2513.4]
  assign _T_3153 = _T_3131 + _T_3132; // @[Bitwise.scala 48:55:@2514.4]
  assign _GEN_621 = {{1'd0}, _T_3130}; // @[Bitwise.scala 48:55:@2515.4]
  assign _T_3154 = _GEN_621 + _T_3153; // @[Bitwise.scala 48:55:@2515.4]
  assign _T_3155 = _T_3152 + _T_3154; // @[Bitwise.scala 48:55:@2516.4]
  assign _T_3156 = _T_3134 + _T_3135; // @[Bitwise.scala 48:55:@2517.4]
  assign _GEN_622 = {{1'd0}, _T_3133}; // @[Bitwise.scala 48:55:@2518.4]
  assign _T_3157 = _GEN_622 + _T_3156; // @[Bitwise.scala 48:55:@2518.4]
  assign _T_3158 = _T_3137 + _T_3138; // @[Bitwise.scala 48:55:@2519.4]
  assign _GEN_623 = {{1'd0}, _T_3136}; // @[Bitwise.scala 48:55:@2520.4]
  assign _T_3159 = _GEN_623 + _T_3158; // @[Bitwise.scala 48:55:@2520.4]
  assign _T_3160 = _T_3157 + _T_3159; // @[Bitwise.scala 48:55:@2521.4]
  assign _T_3161 = _T_3155 + _T_3160; // @[Bitwise.scala 48:55:@2522.4]
  assign _T_3162 = _T_3140 + _T_3141; // @[Bitwise.scala 48:55:@2523.4]
  assign _GEN_624 = {{1'd0}, _T_3139}; // @[Bitwise.scala 48:55:@2524.4]
  assign _T_3163 = _GEN_624 + _T_3162; // @[Bitwise.scala 48:55:@2524.4]
  assign _T_3164 = _T_3143 + _T_3144; // @[Bitwise.scala 48:55:@2525.4]
  assign _GEN_625 = {{1'd0}, _T_3142}; // @[Bitwise.scala 48:55:@2526.4]
  assign _T_3165 = _GEN_625 + _T_3164; // @[Bitwise.scala 48:55:@2526.4]
  assign _T_3166 = _T_3163 + _T_3165; // @[Bitwise.scala 48:55:@2527.4]
  assign _T_3167 = _T_3146 + _T_3147; // @[Bitwise.scala 48:55:@2528.4]
  assign _GEN_626 = {{1'd0}, _T_3145}; // @[Bitwise.scala 48:55:@2529.4]
  assign _T_3168 = _GEN_626 + _T_3167; // @[Bitwise.scala 48:55:@2529.4]
  assign _T_3169 = _T_3149 + _T_3150; // @[Bitwise.scala 48:55:@2530.4]
  assign _GEN_627 = {{1'd0}, _T_3148}; // @[Bitwise.scala 48:55:@2531.4]
  assign _T_3170 = _GEN_627 + _T_3169; // @[Bitwise.scala 48:55:@2531.4]
  assign _T_3171 = _T_3168 + _T_3170; // @[Bitwise.scala 48:55:@2532.4]
  assign _T_3172 = _T_3166 + _T_3171; // @[Bitwise.scala 48:55:@2533.4]
  assign _T_3173 = _T_3161 + _T_3172; // @[Bitwise.scala 48:55:@2534.4]
  assign _T_3237 = _T_1124[24:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2599.4]
  assign _T_3238 = _T_3237[0]; // @[Bitwise.scala 50:65:@2600.4]
  assign _T_3239 = _T_3237[1]; // @[Bitwise.scala 50:65:@2601.4]
  assign _T_3240 = _T_3237[2]; // @[Bitwise.scala 50:65:@2602.4]
  assign _T_3241 = _T_3237[3]; // @[Bitwise.scala 50:65:@2603.4]
  assign _T_3242 = _T_3237[4]; // @[Bitwise.scala 50:65:@2604.4]
  assign _T_3243 = _T_3237[5]; // @[Bitwise.scala 50:65:@2605.4]
  assign _T_3244 = _T_3237[6]; // @[Bitwise.scala 50:65:@2606.4]
  assign _T_3245 = _T_3237[7]; // @[Bitwise.scala 50:65:@2607.4]
  assign _T_3246 = _T_3237[8]; // @[Bitwise.scala 50:65:@2608.4]
  assign _T_3247 = _T_3237[9]; // @[Bitwise.scala 50:65:@2609.4]
  assign _T_3248 = _T_3237[10]; // @[Bitwise.scala 50:65:@2610.4]
  assign _T_3249 = _T_3237[11]; // @[Bitwise.scala 50:65:@2611.4]
  assign _T_3250 = _T_3237[12]; // @[Bitwise.scala 50:65:@2612.4]
  assign _T_3251 = _T_3237[13]; // @[Bitwise.scala 50:65:@2613.4]
  assign _T_3252 = _T_3237[14]; // @[Bitwise.scala 50:65:@2614.4]
  assign _T_3253 = _T_3237[15]; // @[Bitwise.scala 50:65:@2615.4]
  assign _T_3254 = _T_3237[16]; // @[Bitwise.scala 50:65:@2616.4]
  assign _T_3255 = _T_3237[17]; // @[Bitwise.scala 50:65:@2617.4]
  assign _T_3256 = _T_3237[18]; // @[Bitwise.scala 50:65:@2618.4]
  assign _T_3257 = _T_3237[19]; // @[Bitwise.scala 50:65:@2619.4]
  assign _T_3258 = _T_3237[20]; // @[Bitwise.scala 50:65:@2620.4]
  assign _T_3259 = _T_3237[21]; // @[Bitwise.scala 50:65:@2621.4]
  assign _T_3260 = _T_3237[22]; // @[Bitwise.scala 50:65:@2622.4]
  assign _T_3261 = _T_3237[23]; // @[Bitwise.scala 50:65:@2623.4]
  assign _T_3262 = _T_3237[24]; // @[Bitwise.scala 50:65:@2624.4]
  assign _T_3263 = _T_3239 + _T_3240; // @[Bitwise.scala 48:55:@2625.4]
  assign _GEN_628 = {{1'd0}, _T_3238}; // @[Bitwise.scala 48:55:@2626.4]
  assign _T_3264 = _GEN_628 + _T_3263; // @[Bitwise.scala 48:55:@2626.4]
  assign _T_3265 = _T_3242 + _T_3243; // @[Bitwise.scala 48:55:@2627.4]
  assign _GEN_629 = {{1'd0}, _T_3241}; // @[Bitwise.scala 48:55:@2628.4]
  assign _T_3266 = _GEN_629 + _T_3265; // @[Bitwise.scala 48:55:@2628.4]
  assign _T_3267 = _T_3264 + _T_3266; // @[Bitwise.scala 48:55:@2629.4]
  assign _T_3268 = _T_3245 + _T_3246; // @[Bitwise.scala 48:55:@2630.4]
  assign _GEN_630 = {{1'd0}, _T_3244}; // @[Bitwise.scala 48:55:@2631.4]
  assign _T_3269 = _GEN_630 + _T_3268; // @[Bitwise.scala 48:55:@2631.4]
  assign _T_3270 = _T_3248 + _T_3249; // @[Bitwise.scala 48:55:@2632.4]
  assign _GEN_631 = {{1'd0}, _T_3247}; // @[Bitwise.scala 48:55:@2633.4]
  assign _T_3271 = _GEN_631 + _T_3270; // @[Bitwise.scala 48:55:@2633.4]
  assign _T_3272 = _T_3269 + _T_3271; // @[Bitwise.scala 48:55:@2634.4]
  assign _T_3273 = _T_3267 + _T_3272; // @[Bitwise.scala 48:55:@2635.4]
  assign _T_3274 = _T_3251 + _T_3252; // @[Bitwise.scala 48:55:@2636.4]
  assign _GEN_632 = {{1'd0}, _T_3250}; // @[Bitwise.scala 48:55:@2637.4]
  assign _T_3275 = _GEN_632 + _T_3274; // @[Bitwise.scala 48:55:@2637.4]
  assign _T_3276 = _T_3254 + _T_3255; // @[Bitwise.scala 48:55:@2638.4]
  assign _GEN_633 = {{1'd0}, _T_3253}; // @[Bitwise.scala 48:55:@2639.4]
  assign _T_3277 = _GEN_633 + _T_3276; // @[Bitwise.scala 48:55:@2639.4]
  assign _T_3278 = _T_3275 + _T_3277; // @[Bitwise.scala 48:55:@2640.4]
  assign _T_3279 = _T_3257 + _T_3258; // @[Bitwise.scala 48:55:@2641.4]
  assign _GEN_634 = {{1'd0}, _T_3256}; // @[Bitwise.scala 48:55:@2642.4]
  assign _T_3280 = _GEN_634 + _T_3279; // @[Bitwise.scala 48:55:@2642.4]
  assign _T_3281 = _T_3259 + _T_3260; // @[Bitwise.scala 48:55:@2643.4]
  assign _T_3282 = _T_3261 + _T_3262; // @[Bitwise.scala 48:55:@2644.4]
  assign _T_3283 = _T_3281 + _T_3282; // @[Bitwise.scala 48:55:@2645.4]
  assign _T_3284 = _T_3280 + _T_3283; // @[Bitwise.scala 48:55:@2646.4]
  assign _T_3285 = _T_3278 + _T_3284; // @[Bitwise.scala 48:55:@2647.4]
  assign _T_3286 = _T_3273 + _T_3285; // @[Bitwise.scala 48:55:@2648.4]
  assign _T_3350 = _T_1124[25:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2713.4]
  assign _T_3351 = _T_3350[0]; // @[Bitwise.scala 50:65:@2714.4]
  assign _T_3352 = _T_3350[1]; // @[Bitwise.scala 50:65:@2715.4]
  assign _T_3353 = _T_3350[2]; // @[Bitwise.scala 50:65:@2716.4]
  assign _T_3354 = _T_3350[3]; // @[Bitwise.scala 50:65:@2717.4]
  assign _T_3355 = _T_3350[4]; // @[Bitwise.scala 50:65:@2718.4]
  assign _T_3356 = _T_3350[5]; // @[Bitwise.scala 50:65:@2719.4]
  assign _T_3357 = _T_3350[6]; // @[Bitwise.scala 50:65:@2720.4]
  assign _T_3358 = _T_3350[7]; // @[Bitwise.scala 50:65:@2721.4]
  assign _T_3359 = _T_3350[8]; // @[Bitwise.scala 50:65:@2722.4]
  assign _T_3360 = _T_3350[9]; // @[Bitwise.scala 50:65:@2723.4]
  assign _T_3361 = _T_3350[10]; // @[Bitwise.scala 50:65:@2724.4]
  assign _T_3362 = _T_3350[11]; // @[Bitwise.scala 50:65:@2725.4]
  assign _T_3363 = _T_3350[12]; // @[Bitwise.scala 50:65:@2726.4]
  assign _T_3364 = _T_3350[13]; // @[Bitwise.scala 50:65:@2727.4]
  assign _T_3365 = _T_3350[14]; // @[Bitwise.scala 50:65:@2728.4]
  assign _T_3366 = _T_3350[15]; // @[Bitwise.scala 50:65:@2729.4]
  assign _T_3367 = _T_3350[16]; // @[Bitwise.scala 50:65:@2730.4]
  assign _T_3368 = _T_3350[17]; // @[Bitwise.scala 50:65:@2731.4]
  assign _T_3369 = _T_3350[18]; // @[Bitwise.scala 50:65:@2732.4]
  assign _T_3370 = _T_3350[19]; // @[Bitwise.scala 50:65:@2733.4]
  assign _T_3371 = _T_3350[20]; // @[Bitwise.scala 50:65:@2734.4]
  assign _T_3372 = _T_3350[21]; // @[Bitwise.scala 50:65:@2735.4]
  assign _T_3373 = _T_3350[22]; // @[Bitwise.scala 50:65:@2736.4]
  assign _T_3374 = _T_3350[23]; // @[Bitwise.scala 50:65:@2737.4]
  assign _T_3375 = _T_3350[24]; // @[Bitwise.scala 50:65:@2738.4]
  assign _T_3376 = _T_3350[25]; // @[Bitwise.scala 50:65:@2739.4]
  assign _T_3377 = _T_3352 + _T_3353; // @[Bitwise.scala 48:55:@2740.4]
  assign _GEN_635 = {{1'd0}, _T_3351}; // @[Bitwise.scala 48:55:@2741.4]
  assign _T_3378 = _GEN_635 + _T_3377; // @[Bitwise.scala 48:55:@2741.4]
  assign _T_3379 = _T_3355 + _T_3356; // @[Bitwise.scala 48:55:@2742.4]
  assign _GEN_636 = {{1'd0}, _T_3354}; // @[Bitwise.scala 48:55:@2743.4]
  assign _T_3380 = _GEN_636 + _T_3379; // @[Bitwise.scala 48:55:@2743.4]
  assign _T_3381 = _T_3378 + _T_3380; // @[Bitwise.scala 48:55:@2744.4]
  assign _T_3382 = _T_3358 + _T_3359; // @[Bitwise.scala 48:55:@2745.4]
  assign _GEN_637 = {{1'd0}, _T_3357}; // @[Bitwise.scala 48:55:@2746.4]
  assign _T_3383 = _GEN_637 + _T_3382; // @[Bitwise.scala 48:55:@2746.4]
  assign _T_3384 = _T_3360 + _T_3361; // @[Bitwise.scala 48:55:@2747.4]
  assign _T_3385 = _T_3362 + _T_3363; // @[Bitwise.scala 48:55:@2748.4]
  assign _T_3386 = _T_3384 + _T_3385; // @[Bitwise.scala 48:55:@2749.4]
  assign _T_3387 = _T_3383 + _T_3386; // @[Bitwise.scala 48:55:@2750.4]
  assign _T_3388 = _T_3381 + _T_3387; // @[Bitwise.scala 48:55:@2751.4]
  assign _T_3389 = _T_3365 + _T_3366; // @[Bitwise.scala 48:55:@2752.4]
  assign _GEN_638 = {{1'd0}, _T_3364}; // @[Bitwise.scala 48:55:@2753.4]
  assign _T_3390 = _GEN_638 + _T_3389; // @[Bitwise.scala 48:55:@2753.4]
  assign _T_3391 = _T_3368 + _T_3369; // @[Bitwise.scala 48:55:@2754.4]
  assign _GEN_639 = {{1'd0}, _T_3367}; // @[Bitwise.scala 48:55:@2755.4]
  assign _T_3392 = _GEN_639 + _T_3391; // @[Bitwise.scala 48:55:@2755.4]
  assign _T_3393 = _T_3390 + _T_3392; // @[Bitwise.scala 48:55:@2756.4]
  assign _T_3394 = _T_3371 + _T_3372; // @[Bitwise.scala 48:55:@2757.4]
  assign _GEN_640 = {{1'd0}, _T_3370}; // @[Bitwise.scala 48:55:@2758.4]
  assign _T_3395 = _GEN_640 + _T_3394; // @[Bitwise.scala 48:55:@2758.4]
  assign _T_3396 = _T_3373 + _T_3374; // @[Bitwise.scala 48:55:@2759.4]
  assign _T_3397 = _T_3375 + _T_3376; // @[Bitwise.scala 48:55:@2760.4]
  assign _T_3398 = _T_3396 + _T_3397; // @[Bitwise.scala 48:55:@2761.4]
  assign _T_3399 = _T_3395 + _T_3398; // @[Bitwise.scala 48:55:@2762.4]
  assign _T_3400 = _T_3393 + _T_3399; // @[Bitwise.scala 48:55:@2763.4]
  assign _T_3401 = _T_3388 + _T_3400; // @[Bitwise.scala 48:55:@2764.4]
  assign _T_3465 = _T_1124[26:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2829.4]
  assign _T_3466 = _T_3465[0]; // @[Bitwise.scala 50:65:@2830.4]
  assign _T_3467 = _T_3465[1]; // @[Bitwise.scala 50:65:@2831.4]
  assign _T_3468 = _T_3465[2]; // @[Bitwise.scala 50:65:@2832.4]
  assign _T_3469 = _T_3465[3]; // @[Bitwise.scala 50:65:@2833.4]
  assign _T_3470 = _T_3465[4]; // @[Bitwise.scala 50:65:@2834.4]
  assign _T_3471 = _T_3465[5]; // @[Bitwise.scala 50:65:@2835.4]
  assign _T_3472 = _T_3465[6]; // @[Bitwise.scala 50:65:@2836.4]
  assign _T_3473 = _T_3465[7]; // @[Bitwise.scala 50:65:@2837.4]
  assign _T_3474 = _T_3465[8]; // @[Bitwise.scala 50:65:@2838.4]
  assign _T_3475 = _T_3465[9]; // @[Bitwise.scala 50:65:@2839.4]
  assign _T_3476 = _T_3465[10]; // @[Bitwise.scala 50:65:@2840.4]
  assign _T_3477 = _T_3465[11]; // @[Bitwise.scala 50:65:@2841.4]
  assign _T_3478 = _T_3465[12]; // @[Bitwise.scala 50:65:@2842.4]
  assign _T_3479 = _T_3465[13]; // @[Bitwise.scala 50:65:@2843.4]
  assign _T_3480 = _T_3465[14]; // @[Bitwise.scala 50:65:@2844.4]
  assign _T_3481 = _T_3465[15]; // @[Bitwise.scala 50:65:@2845.4]
  assign _T_3482 = _T_3465[16]; // @[Bitwise.scala 50:65:@2846.4]
  assign _T_3483 = _T_3465[17]; // @[Bitwise.scala 50:65:@2847.4]
  assign _T_3484 = _T_3465[18]; // @[Bitwise.scala 50:65:@2848.4]
  assign _T_3485 = _T_3465[19]; // @[Bitwise.scala 50:65:@2849.4]
  assign _T_3486 = _T_3465[20]; // @[Bitwise.scala 50:65:@2850.4]
  assign _T_3487 = _T_3465[21]; // @[Bitwise.scala 50:65:@2851.4]
  assign _T_3488 = _T_3465[22]; // @[Bitwise.scala 50:65:@2852.4]
  assign _T_3489 = _T_3465[23]; // @[Bitwise.scala 50:65:@2853.4]
  assign _T_3490 = _T_3465[24]; // @[Bitwise.scala 50:65:@2854.4]
  assign _T_3491 = _T_3465[25]; // @[Bitwise.scala 50:65:@2855.4]
  assign _T_3492 = _T_3465[26]; // @[Bitwise.scala 50:65:@2856.4]
  assign _T_3493 = _T_3467 + _T_3468; // @[Bitwise.scala 48:55:@2857.4]
  assign _GEN_641 = {{1'd0}, _T_3466}; // @[Bitwise.scala 48:55:@2858.4]
  assign _T_3494 = _GEN_641 + _T_3493; // @[Bitwise.scala 48:55:@2858.4]
  assign _T_3495 = _T_3470 + _T_3471; // @[Bitwise.scala 48:55:@2859.4]
  assign _GEN_642 = {{1'd0}, _T_3469}; // @[Bitwise.scala 48:55:@2860.4]
  assign _T_3496 = _GEN_642 + _T_3495; // @[Bitwise.scala 48:55:@2860.4]
  assign _T_3497 = _T_3494 + _T_3496; // @[Bitwise.scala 48:55:@2861.4]
  assign _T_3498 = _T_3473 + _T_3474; // @[Bitwise.scala 48:55:@2862.4]
  assign _GEN_643 = {{1'd0}, _T_3472}; // @[Bitwise.scala 48:55:@2863.4]
  assign _T_3499 = _GEN_643 + _T_3498; // @[Bitwise.scala 48:55:@2863.4]
  assign _T_3500 = _T_3475 + _T_3476; // @[Bitwise.scala 48:55:@2864.4]
  assign _T_3501 = _T_3477 + _T_3478; // @[Bitwise.scala 48:55:@2865.4]
  assign _T_3502 = _T_3500 + _T_3501; // @[Bitwise.scala 48:55:@2866.4]
  assign _T_3503 = _T_3499 + _T_3502; // @[Bitwise.scala 48:55:@2867.4]
  assign _T_3504 = _T_3497 + _T_3503; // @[Bitwise.scala 48:55:@2868.4]
  assign _T_3505 = _T_3480 + _T_3481; // @[Bitwise.scala 48:55:@2869.4]
  assign _GEN_644 = {{1'd0}, _T_3479}; // @[Bitwise.scala 48:55:@2870.4]
  assign _T_3506 = _GEN_644 + _T_3505; // @[Bitwise.scala 48:55:@2870.4]
  assign _T_3507 = _T_3482 + _T_3483; // @[Bitwise.scala 48:55:@2871.4]
  assign _T_3508 = _T_3484 + _T_3485; // @[Bitwise.scala 48:55:@2872.4]
  assign _T_3509 = _T_3507 + _T_3508; // @[Bitwise.scala 48:55:@2873.4]
  assign _T_3510 = _T_3506 + _T_3509; // @[Bitwise.scala 48:55:@2874.4]
  assign _T_3511 = _T_3487 + _T_3488; // @[Bitwise.scala 48:55:@2875.4]
  assign _GEN_645 = {{1'd0}, _T_3486}; // @[Bitwise.scala 48:55:@2876.4]
  assign _T_3512 = _GEN_645 + _T_3511; // @[Bitwise.scala 48:55:@2876.4]
  assign _T_3513 = _T_3489 + _T_3490; // @[Bitwise.scala 48:55:@2877.4]
  assign _T_3514 = _T_3491 + _T_3492; // @[Bitwise.scala 48:55:@2878.4]
  assign _T_3515 = _T_3513 + _T_3514; // @[Bitwise.scala 48:55:@2879.4]
  assign _T_3516 = _T_3512 + _T_3515; // @[Bitwise.scala 48:55:@2880.4]
  assign _T_3517 = _T_3510 + _T_3516; // @[Bitwise.scala 48:55:@2881.4]
  assign _T_3518 = _T_3504 + _T_3517; // @[Bitwise.scala 48:55:@2882.4]
  assign _T_3582 = _T_1124[27:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@2947.4]
  assign _T_3583 = _T_3582[0]; // @[Bitwise.scala 50:65:@2948.4]
  assign _T_3584 = _T_3582[1]; // @[Bitwise.scala 50:65:@2949.4]
  assign _T_3585 = _T_3582[2]; // @[Bitwise.scala 50:65:@2950.4]
  assign _T_3586 = _T_3582[3]; // @[Bitwise.scala 50:65:@2951.4]
  assign _T_3587 = _T_3582[4]; // @[Bitwise.scala 50:65:@2952.4]
  assign _T_3588 = _T_3582[5]; // @[Bitwise.scala 50:65:@2953.4]
  assign _T_3589 = _T_3582[6]; // @[Bitwise.scala 50:65:@2954.4]
  assign _T_3590 = _T_3582[7]; // @[Bitwise.scala 50:65:@2955.4]
  assign _T_3591 = _T_3582[8]; // @[Bitwise.scala 50:65:@2956.4]
  assign _T_3592 = _T_3582[9]; // @[Bitwise.scala 50:65:@2957.4]
  assign _T_3593 = _T_3582[10]; // @[Bitwise.scala 50:65:@2958.4]
  assign _T_3594 = _T_3582[11]; // @[Bitwise.scala 50:65:@2959.4]
  assign _T_3595 = _T_3582[12]; // @[Bitwise.scala 50:65:@2960.4]
  assign _T_3596 = _T_3582[13]; // @[Bitwise.scala 50:65:@2961.4]
  assign _T_3597 = _T_3582[14]; // @[Bitwise.scala 50:65:@2962.4]
  assign _T_3598 = _T_3582[15]; // @[Bitwise.scala 50:65:@2963.4]
  assign _T_3599 = _T_3582[16]; // @[Bitwise.scala 50:65:@2964.4]
  assign _T_3600 = _T_3582[17]; // @[Bitwise.scala 50:65:@2965.4]
  assign _T_3601 = _T_3582[18]; // @[Bitwise.scala 50:65:@2966.4]
  assign _T_3602 = _T_3582[19]; // @[Bitwise.scala 50:65:@2967.4]
  assign _T_3603 = _T_3582[20]; // @[Bitwise.scala 50:65:@2968.4]
  assign _T_3604 = _T_3582[21]; // @[Bitwise.scala 50:65:@2969.4]
  assign _T_3605 = _T_3582[22]; // @[Bitwise.scala 50:65:@2970.4]
  assign _T_3606 = _T_3582[23]; // @[Bitwise.scala 50:65:@2971.4]
  assign _T_3607 = _T_3582[24]; // @[Bitwise.scala 50:65:@2972.4]
  assign _T_3608 = _T_3582[25]; // @[Bitwise.scala 50:65:@2973.4]
  assign _T_3609 = _T_3582[26]; // @[Bitwise.scala 50:65:@2974.4]
  assign _T_3610 = _T_3582[27]; // @[Bitwise.scala 50:65:@2975.4]
  assign _T_3611 = _T_3584 + _T_3585; // @[Bitwise.scala 48:55:@2976.4]
  assign _GEN_646 = {{1'd0}, _T_3583}; // @[Bitwise.scala 48:55:@2977.4]
  assign _T_3612 = _GEN_646 + _T_3611; // @[Bitwise.scala 48:55:@2977.4]
  assign _T_3613 = _T_3586 + _T_3587; // @[Bitwise.scala 48:55:@2978.4]
  assign _T_3614 = _T_3588 + _T_3589; // @[Bitwise.scala 48:55:@2979.4]
  assign _T_3615 = _T_3613 + _T_3614; // @[Bitwise.scala 48:55:@2980.4]
  assign _T_3616 = _T_3612 + _T_3615; // @[Bitwise.scala 48:55:@2981.4]
  assign _T_3617 = _T_3591 + _T_3592; // @[Bitwise.scala 48:55:@2982.4]
  assign _GEN_647 = {{1'd0}, _T_3590}; // @[Bitwise.scala 48:55:@2983.4]
  assign _T_3618 = _GEN_647 + _T_3617; // @[Bitwise.scala 48:55:@2983.4]
  assign _T_3619 = _T_3593 + _T_3594; // @[Bitwise.scala 48:55:@2984.4]
  assign _T_3620 = _T_3595 + _T_3596; // @[Bitwise.scala 48:55:@2985.4]
  assign _T_3621 = _T_3619 + _T_3620; // @[Bitwise.scala 48:55:@2986.4]
  assign _T_3622 = _T_3618 + _T_3621; // @[Bitwise.scala 48:55:@2987.4]
  assign _T_3623 = _T_3616 + _T_3622; // @[Bitwise.scala 48:55:@2988.4]
  assign _T_3624 = _T_3598 + _T_3599; // @[Bitwise.scala 48:55:@2989.4]
  assign _GEN_648 = {{1'd0}, _T_3597}; // @[Bitwise.scala 48:55:@2990.4]
  assign _T_3625 = _GEN_648 + _T_3624; // @[Bitwise.scala 48:55:@2990.4]
  assign _T_3626 = _T_3600 + _T_3601; // @[Bitwise.scala 48:55:@2991.4]
  assign _T_3627 = _T_3602 + _T_3603; // @[Bitwise.scala 48:55:@2992.4]
  assign _T_3628 = _T_3626 + _T_3627; // @[Bitwise.scala 48:55:@2993.4]
  assign _T_3629 = _T_3625 + _T_3628; // @[Bitwise.scala 48:55:@2994.4]
  assign _T_3630 = _T_3605 + _T_3606; // @[Bitwise.scala 48:55:@2995.4]
  assign _GEN_649 = {{1'd0}, _T_3604}; // @[Bitwise.scala 48:55:@2996.4]
  assign _T_3631 = _GEN_649 + _T_3630; // @[Bitwise.scala 48:55:@2996.4]
  assign _T_3632 = _T_3607 + _T_3608; // @[Bitwise.scala 48:55:@2997.4]
  assign _T_3633 = _T_3609 + _T_3610; // @[Bitwise.scala 48:55:@2998.4]
  assign _T_3634 = _T_3632 + _T_3633; // @[Bitwise.scala 48:55:@2999.4]
  assign _T_3635 = _T_3631 + _T_3634; // @[Bitwise.scala 48:55:@3000.4]
  assign _T_3636 = _T_3629 + _T_3635; // @[Bitwise.scala 48:55:@3001.4]
  assign _T_3637 = _T_3623 + _T_3636; // @[Bitwise.scala 48:55:@3002.4]
  assign _T_3701 = _T_1124[28:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3067.4]
  assign _T_3702 = _T_3701[0]; // @[Bitwise.scala 50:65:@3068.4]
  assign _T_3703 = _T_3701[1]; // @[Bitwise.scala 50:65:@3069.4]
  assign _T_3704 = _T_3701[2]; // @[Bitwise.scala 50:65:@3070.4]
  assign _T_3705 = _T_3701[3]; // @[Bitwise.scala 50:65:@3071.4]
  assign _T_3706 = _T_3701[4]; // @[Bitwise.scala 50:65:@3072.4]
  assign _T_3707 = _T_3701[5]; // @[Bitwise.scala 50:65:@3073.4]
  assign _T_3708 = _T_3701[6]; // @[Bitwise.scala 50:65:@3074.4]
  assign _T_3709 = _T_3701[7]; // @[Bitwise.scala 50:65:@3075.4]
  assign _T_3710 = _T_3701[8]; // @[Bitwise.scala 50:65:@3076.4]
  assign _T_3711 = _T_3701[9]; // @[Bitwise.scala 50:65:@3077.4]
  assign _T_3712 = _T_3701[10]; // @[Bitwise.scala 50:65:@3078.4]
  assign _T_3713 = _T_3701[11]; // @[Bitwise.scala 50:65:@3079.4]
  assign _T_3714 = _T_3701[12]; // @[Bitwise.scala 50:65:@3080.4]
  assign _T_3715 = _T_3701[13]; // @[Bitwise.scala 50:65:@3081.4]
  assign _T_3716 = _T_3701[14]; // @[Bitwise.scala 50:65:@3082.4]
  assign _T_3717 = _T_3701[15]; // @[Bitwise.scala 50:65:@3083.4]
  assign _T_3718 = _T_3701[16]; // @[Bitwise.scala 50:65:@3084.4]
  assign _T_3719 = _T_3701[17]; // @[Bitwise.scala 50:65:@3085.4]
  assign _T_3720 = _T_3701[18]; // @[Bitwise.scala 50:65:@3086.4]
  assign _T_3721 = _T_3701[19]; // @[Bitwise.scala 50:65:@3087.4]
  assign _T_3722 = _T_3701[20]; // @[Bitwise.scala 50:65:@3088.4]
  assign _T_3723 = _T_3701[21]; // @[Bitwise.scala 50:65:@3089.4]
  assign _T_3724 = _T_3701[22]; // @[Bitwise.scala 50:65:@3090.4]
  assign _T_3725 = _T_3701[23]; // @[Bitwise.scala 50:65:@3091.4]
  assign _T_3726 = _T_3701[24]; // @[Bitwise.scala 50:65:@3092.4]
  assign _T_3727 = _T_3701[25]; // @[Bitwise.scala 50:65:@3093.4]
  assign _T_3728 = _T_3701[26]; // @[Bitwise.scala 50:65:@3094.4]
  assign _T_3729 = _T_3701[27]; // @[Bitwise.scala 50:65:@3095.4]
  assign _T_3730 = _T_3701[28]; // @[Bitwise.scala 50:65:@3096.4]
  assign _T_3731 = _T_3703 + _T_3704; // @[Bitwise.scala 48:55:@3097.4]
  assign _GEN_650 = {{1'd0}, _T_3702}; // @[Bitwise.scala 48:55:@3098.4]
  assign _T_3732 = _GEN_650 + _T_3731; // @[Bitwise.scala 48:55:@3098.4]
  assign _T_3733 = _T_3705 + _T_3706; // @[Bitwise.scala 48:55:@3099.4]
  assign _T_3734 = _T_3707 + _T_3708; // @[Bitwise.scala 48:55:@3100.4]
  assign _T_3735 = _T_3733 + _T_3734; // @[Bitwise.scala 48:55:@3101.4]
  assign _T_3736 = _T_3732 + _T_3735; // @[Bitwise.scala 48:55:@3102.4]
  assign _T_3737 = _T_3710 + _T_3711; // @[Bitwise.scala 48:55:@3103.4]
  assign _GEN_651 = {{1'd0}, _T_3709}; // @[Bitwise.scala 48:55:@3104.4]
  assign _T_3738 = _GEN_651 + _T_3737; // @[Bitwise.scala 48:55:@3104.4]
  assign _T_3739 = _T_3712 + _T_3713; // @[Bitwise.scala 48:55:@3105.4]
  assign _T_3740 = _T_3714 + _T_3715; // @[Bitwise.scala 48:55:@3106.4]
  assign _T_3741 = _T_3739 + _T_3740; // @[Bitwise.scala 48:55:@3107.4]
  assign _T_3742 = _T_3738 + _T_3741; // @[Bitwise.scala 48:55:@3108.4]
  assign _T_3743 = _T_3736 + _T_3742; // @[Bitwise.scala 48:55:@3109.4]
  assign _T_3744 = _T_3717 + _T_3718; // @[Bitwise.scala 48:55:@3110.4]
  assign _GEN_652 = {{1'd0}, _T_3716}; // @[Bitwise.scala 48:55:@3111.4]
  assign _T_3745 = _GEN_652 + _T_3744; // @[Bitwise.scala 48:55:@3111.4]
  assign _T_3746 = _T_3719 + _T_3720; // @[Bitwise.scala 48:55:@3112.4]
  assign _T_3747 = _T_3721 + _T_3722; // @[Bitwise.scala 48:55:@3113.4]
  assign _T_3748 = _T_3746 + _T_3747; // @[Bitwise.scala 48:55:@3114.4]
  assign _T_3749 = _T_3745 + _T_3748; // @[Bitwise.scala 48:55:@3115.4]
  assign _T_3750 = _T_3723 + _T_3724; // @[Bitwise.scala 48:55:@3116.4]
  assign _T_3751 = _T_3725 + _T_3726; // @[Bitwise.scala 48:55:@3117.4]
  assign _T_3752 = _T_3750 + _T_3751; // @[Bitwise.scala 48:55:@3118.4]
  assign _T_3753 = _T_3727 + _T_3728; // @[Bitwise.scala 48:55:@3119.4]
  assign _T_3754 = _T_3729 + _T_3730; // @[Bitwise.scala 48:55:@3120.4]
  assign _T_3755 = _T_3753 + _T_3754; // @[Bitwise.scala 48:55:@3121.4]
  assign _T_3756 = _T_3752 + _T_3755; // @[Bitwise.scala 48:55:@3122.4]
  assign _T_3757 = _T_3749 + _T_3756; // @[Bitwise.scala 48:55:@3123.4]
  assign _T_3758 = _T_3743 + _T_3757; // @[Bitwise.scala 48:55:@3124.4]
  assign _T_3822 = _T_1124[29:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3189.4]
  assign _T_3823 = _T_3822[0]; // @[Bitwise.scala 50:65:@3190.4]
  assign _T_3824 = _T_3822[1]; // @[Bitwise.scala 50:65:@3191.4]
  assign _T_3825 = _T_3822[2]; // @[Bitwise.scala 50:65:@3192.4]
  assign _T_3826 = _T_3822[3]; // @[Bitwise.scala 50:65:@3193.4]
  assign _T_3827 = _T_3822[4]; // @[Bitwise.scala 50:65:@3194.4]
  assign _T_3828 = _T_3822[5]; // @[Bitwise.scala 50:65:@3195.4]
  assign _T_3829 = _T_3822[6]; // @[Bitwise.scala 50:65:@3196.4]
  assign _T_3830 = _T_3822[7]; // @[Bitwise.scala 50:65:@3197.4]
  assign _T_3831 = _T_3822[8]; // @[Bitwise.scala 50:65:@3198.4]
  assign _T_3832 = _T_3822[9]; // @[Bitwise.scala 50:65:@3199.4]
  assign _T_3833 = _T_3822[10]; // @[Bitwise.scala 50:65:@3200.4]
  assign _T_3834 = _T_3822[11]; // @[Bitwise.scala 50:65:@3201.4]
  assign _T_3835 = _T_3822[12]; // @[Bitwise.scala 50:65:@3202.4]
  assign _T_3836 = _T_3822[13]; // @[Bitwise.scala 50:65:@3203.4]
  assign _T_3837 = _T_3822[14]; // @[Bitwise.scala 50:65:@3204.4]
  assign _T_3838 = _T_3822[15]; // @[Bitwise.scala 50:65:@3205.4]
  assign _T_3839 = _T_3822[16]; // @[Bitwise.scala 50:65:@3206.4]
  assign _T_3840 = _T_3822[17]; // @[Bitwise.scala 50:65:@3207.4]
  assign _T_3841 = _T_3822[18]; // @[Bitwise.scala 50:65:@3208.4]
  assign _T_3842 = _T_3822[19]; // @[Bitwise.scala 50:65:@3209.4]
  assign _T_3843 = _T_3822[20]; // @[Bitwise.scala 50:65:@3210.4]
  assign _T_3844 = _T_3822[21]; // @[Bitwise.scala 50:65:@3211.4]
  assign _T_3845 = _T_3822[22]; // @[Bitwise.scala 50:65:@3212.4]
  assign _T_3846 = _T_3822[23]; // @[Bitwise.scala 50:65:@3213.4]
  assign _T_3847 = _T_3822[24]; // @[Bitwise.scala 50:65:@3214.4]
  assign _T_3848 = _T_3822[25]; // @[Bitwise.scala 50:65:@3215.4]
  assign _T_3849 = _T_3822[26]; // @[Bitwise.scala 50:65:@3216.4]
  assign _T_3850 = _T_3822[27]; // @[Bitwise.scala 50:65:@3217.4]
  assign _T_3851 = _T_3822[28]; // @[Bitwise.scala 50:65:@3218.4]
  assign _T_3852 = _T_3822[29]; // @[Bitwise.scala 50:65:@3219.4]
  assign _T_3853 = _T_3824 + _T_3825; // @[Bitwise.scala 48:55:@3220.4]
  assign _GEN_653 = {{1'd0}, _T_3823}; // @[Bitwise.scala 48:55:@3221.4]
  assign _T_3854 = _GEN_653 + _T_3853; // @[Bitwise.scala 48:55:@3221.4]
  assign _T_3855 = _T_3826 + _T_3827; // @[Bitwise.scala 48:55:@3222.4]
  assign _T_3856 = _T_3828 + _T_3829; // @[Bitwise.scala 48:55:@3223.4]
  assign _T_3857 = _T_3855 + _T_3856; // @[Bitwise.scala 48:55:@3224.4]
  assign _T_3858 = _T_3854 + _T_3857; // @[Bitwise.scala 48:55:@3225.4]
  assign _T_3859 = _T_3830 + _T_3831; // @[Bitwise.scala 48:55:@3226.4]
  assign _T_3860 = _T_3832 + _T_3833; // @[Bitwise.scala 48:55:@3227.4]
  assign _T_3861 = _T_3859 + _T_3860; // @[Bitwise.scala 48:55:@3228.4]
  assign _T_3862 = _T_3834 + _T_3835; // @[Bitwise.scala 48:55:@3229.4]
  assign _T_3863 = _T_3836 + _T_3837; // @[Bitwise.scala 48:55:@3230.4]
  assign _T_3864 = _T_3862 + _T_3863; // @[Bitwise.scala 48:55:@3231.4]
  assign _T_3865 = _T_3861 + _T_3864; // @[Bitwise.scala 48:55:@3232.4]
  assign _T_3866 = _T_3858 + _T_3865; // @[Bitwise.scala 48:55:@3233.4]
  assign _T_3867 = _T_3839 + _T_3840; // @[Bitwise.scala 48:55:@3234.4]
  assign _GEN_654 = {{1'd0}, _T_3838}; // @[Bitwise.scala 48:55:@3235.4]
  assign _T_3868 = _GEN_654 + _T_3867; // @[Bitwise.scala 48:55:@3235.4]
  assign _T_3869 = _T_3841 + _T_3842; // @[Bitwise.scala 48:55:@3236.4]
  assign _T_3870 = _T_3843 + _T_3844; // @[Bitwise.scala 48:55:@3237.4]
  assign _T_3871 = _T_3869 + _T_3870; // @[Bitwise.scala 48:55:@3238.4]
  assign _T_3872 = _T_3868 + _T_3871; // @[Bitwise.scala 48:55:@3239.4]
  assign _T_3873 = _T_3845 + _T_3846; // @[Bitwise.scala 48:55:@3240.4]
  assign _T_3874 = _T_3847 + _T_3848; // @[Bitwise.scala 48:55:@3241.4]
  assign _T_3875 = _T_3873 + _T_3874; // @[Bitwise.scala 48:55:@3242.4]
  assign _T_3876 = _T_3849 + _T_3850; // @[Bitwise.scala 48:55:@3243.4]
  assign _T_3877 = _T_3851 + _T_3852; // @[Bitwise.scala 48:55:@3244.4]
  assign _T_3878 = _T_3876 + _T_3877; // @[Bitwise.scala 48:55:@3245.4]
  assign _T_3879 = _T_3875 + _T_3878; // @[Bitwise.scala 48:55:@3246.4]
  assign _T_3880 = _T_3872 + _T_3879; // @[Bitwise.scala 48:55:@3247.4]
  assign _T_3881 = _T_3866 + _T_3880; // @[Bitwise.scala 48:55:@3248.4]
  assign _T_3945 = _T_1124[30:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3313.4]
  assign _T_3946 = _T_3945[0]; // @[Bitwise.scala 50:65:@3314.4]
  assign _T_3947 = _T_3945[1]; // @[Bitwise.scala 50:65:@3315.4]
  assign _T_3948 = _T_3945[2]; // @[Bitwise.scala 50:65:@3316.4]
  assign _T_3949 = _T_3945[3]; // @[Bitwise.scala 50:65:@3317.4]
  assign _T_3950 = _T_3945[4]; // @[Bitwise.scala 50:65:@3318.4]
  assign _T_3951 = _T_3945[5]; // @[Bitwise.scala 50:65:@3319.4]
  assign _T_3952 = _T_3945[6]; // @[Bitwise.scala 50:65:@3320.4]
  assign _T_3953 = _T_3945[7]; // @[Bitwise.scala 50:65:@3321.4]
  assign _T_3954 = _T_3945[8]; // @[Bitwise.scala 50:65:@3322.4]
  assign _T_3955 = _T_3945[9]; // @[Bitwise.scala 50:65:@3323.4]
  assign _T_3956 = _T_3945[10]; // @[Bitwise.scala 50:65:@3324.4]
  assign _T_3957 = _T_3945[11]; // @[Bitwise.scala 50:65:@3325.4]
  assign _T_3958 = _T_3945[12]; // @[Bitwise.scala 50:65:@3326.4]
  assign _T_3959 = _T_3945[13]; // @[Bitwise.scala 50:65:@3327.4]
  assign _T_3960 = _T_3945[14]; // @[Bitwise.scala 50:65:@3328.4]
  assign _T_3961 = _T_3945[15]; // @[Bitwise.scala 50:65:@3329.4]
  assign _T_3962 = _T_3945[16]; // @[Bitwise.scala 50:65:@3330.4]
  assign _T_3963 = _T_3945[17]; // @[Bitwise.scala 50:65:@3331.4]
  assign _T_3964 = _T_3945[18]; // @[Bitwise.scala 50:65:@3332.4]
  assign _T_3965 = _T_3945[19]; // @[Bitwise.scala 50:65:@3333.4]
  assign _T_3966 = _T_3945[20]; // @[Bitwise.scala 50:65:@3334.4]
  assign _T_3967 = _T_3945[21]; // @[Bitwise.scala 50:65:@3335.4]
  assign _T_3968 = _T_3945[22]; // @[Bitwise.scala 50:65:@3336.4]
  assign _T_3969 = _T_3945[23]; // @[Bitwise.scala 50:65:@3337.4]
  assign _T_3970 = _T_3945[24]; // @[Bitwise.scala 50:65:@3338.4]
  assign _T_3971 = _T_3945[25]; // @[Bitwise.scala 50:65:@3339.4]
  assign _T_3972 = _T_3945[26]; // @[Bitwise.scala 50:65:@3340.4]
  assign _T_3973 = _T_3945[27]; // @[Bitwise.scala 50:65:@3341.4]
  assign _T_3974 = _T_3945[28]; // @[Bitwise.scala 50:65:@3342.4]
  assign _T_3975 = _T_3945[29]; // @[Bitwise.scala 50:65:@3343.4]
  assign _T_3976 = _T_3945[30]; // @[Bitwise.scala 50:65:@3344.4]
  assign _T_3977 = _T_3947 + _T_3948; // @[Bitwise.scala 48:55:@3345.4]
  assign _GEN_655 = {{1'd0}, _T_3946}; // @[Bitwise.scala 48:55:@3346.4]
  assign _T_3978 = _GEN_655 + _T_3977; // @[Bitwise.scala 48:55:@3346.4]
  assign _T_3979 = _T_3949 + _T_3950; // @[Bitwise.scala 48:55:@3347.4]
  assign _T_3980 = _T_3951 + _T_3952; // @[Bitwise.scala 48:55:@3348.4]
  assign _T_3981 = _T_3979 + _T_3980; // @[Bitwise.scala 48:55:@3349.4]
  assign _T_3982 = _T_3978 + _T_3981; // @[Bitwise.scala 48:55:@3350.4]
  assign _T_3983 = _T_3953 + _T_3954; // @[Bitwise.scala 48:55:@3351.4]
  assign _T_3984 = _T_3955 + _T_3956; // @[Bitwise.scala 48:55:@3352.4]
  assign _T_3985 = _T_3983 + _T_3984; // @[Bitwise.scala 48:55:@3353.4]
  assign _T_3986 = _T_3957 + _T_3958; // @[Bitwise.scala 48:55:@3354.4]
  assign _T_3987 = _T_3959 + _T_3960; // @[Bitwise.scala 48:55:@3355.4]
  assign _T_3988 = _T_3986 + _T_3987; // @[Bitwise.scala 48:55:@3356.4]
  assign _T_3989 = _T_3985 + _T_3988; // @[Bitwise.scala 48:55:@3357.4]
  assign _T_3990 = _T_3982 + _T_3989; // @[Bitwise.scala 48:55:@3358.4]
  assign _T_3991 = _T_3961 + _T_3962; // @[Bitwise.scala 48:55:@3359.4]
  assign _T_3992 = _T_3963 + _T_3964; // @[Bitwise.scala 48:55:@3360.4]
  assign _T_3993 = _T_3991 + _T_3992; // @[Bitwise.scala 48:55:@3361.4]
  assign _T_3994 = _T_3965 + _T_3966; // @[Bitwise.scala 48:55:@3362.4]
  assign _T_3995 = _T_3967 + _T_3968; // @[Bitwise.scala 48:55:@3363.4]
  assign _T_3996 = _T_3994 + _T_3995; // @[Bitwise.scala 48:55:@3364.4]
  assign _T_3997 = _T_3993 + _T_3996; // @[Bitwise.scala 48:55:@3365.4]
  assign _T_3998 = _T_3969 + _T_3970; // @[Bitwise.scala 48:55:@3366.4]
  assign _T_3999 = _T_3971 + _T_3972; // @[Bitwise.scala 48:55:@3367.4]
  assign _T_4000 = _T_3998 + _T_3999; // @[Bitwise.scala 48:55:@3368.4]
  assign _T_4001 = _T_3973 + _T_3974; // @[Bitwise.scala 48:55:@3369.4]
  assign _T_4002 = _T_3975 + _T_3976; // @[Bitwise.scala 48:55:@3370.4]
  assign _T_4003 = _T_4001 + _T_4002; // @[Bitwise.scala 48:55:@3371.4]
  assign _T_4004 = _T_4000 + _T_4003; // @[Bitwise.scala 48:55:@3372.4]
  assign _T_4005 = _T_3997 + _T_4004; // @[Bitwise.scala 48:55:@3373.4]
  assign _T_4006 = _T_3990 + _T_4005; // @[Bitwise.scala 48:55:@3374.4]
  assign _T_4070 = _T_1124[31:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3439.4]
  assign _T_4071 = _T_4070[0]; // @[Bitwise.scala 50:65:@3440.4]
  assign _T_4072 = _T_4070[1]; // @[Bitwise.scala 50:65:@3441.4]
  assign _T_4073 = _T_4070[2]; // @[Bitwise.scala 50:65:@3442.4]
  assign _T_4074 = _T_4070[3]; // @[Bitwise.scala 50:65:@3443.4]
  assign _T_4075 = _T_4070[4]; // @[Bitwise.scala 50:65:@3444.4]
  assign _T_4076 = _T_4070[5]; // @[Bitwise.scala 50:65:@3445.4]
  assign _T_4077 = _T_4070[6]; // @[Bitwise.scala 50:65:@3446.4]
  assign _T_4078 = _T_4070[7]; // @[Bitwise.scala 50:65:@3447.4]
  assign _T_4079 = _T_4070[8]; // @[Bitwise.scala 50:65:@3448.4]
  assign _T_4080 = _T_4070[9]; // @[Bitwise.scala 50:65:@3449.4]
  assign _T_4081 = _T_4070[10]; // @[Bitwise.scala 50:65:@3450.4]
  assign _T_4082 = _T_4070[11]; // @[Bitwise.scala 50:65:@3451.4]
  assign _T_4083 = _T_4070[12]; // @[Bitwise.scala 50:65:@3452.4]
  assign _T_4084 = _T_4070[13]; // @[Bitwise.scala 50:65:@3453.4]
  assign _T_4085 = _T_4070[14]; // @[Bitwise.scala 50:65:@3454.4]
  assign _T_4086 = _T_4070[15]; // @[Bitwise.scala 50:65:@3455.4]
  assign _T_4087 = _T_4070[16]; // @[Bitwise.scala 50:65:@3456.4]
  assign _T_4088 = _T_4070[17]; // @[Bitwise.scala 50:65:@3457.4]
  assign _T_4089 = _T_4070[18]; // @[Bitwise.scala 50:65:@3458.4]
  assign _T_4090 = _T_4070[19]; // @[Bitwise.scala 50:65:@3459.4]
  assign _T_4091 = _T_4070[20]; // @[Bitwise.scala 50:65:@3460.4]
  assign _T_4092 = _T_4070[21]; // @[Bitwise.scala 50:65:@3461.4]
  assign _T_4093 = _T_4070[22]; // @[Bitwise.scala 50:65:@3462.4]
  assign _T_4094 = _T_4070[23]; // @[Bitwise.scala 50:65:@3463.4]
  assign _T_4095 = _T_4070[24]; // @[Bitwise.scala 50:65:@3464.4]
  assign _T_4096 = _T_4070[25]; // @[Bitwise.scala 50:65:@3465.4]
  assign _T_4097 = _T_4070[26]; // @[Bitwise.scala 50:65:@3466.4]
  assign _T_4098 = _T_4070[27]; // @[Bitwise.scala 50:65:@3467.4]
  assign _T_4099 = _T_4070[28]; // @[Bitwise.scala 50:65:@3468.4]
  assign _T_4100 = _T_4070[29]; // @[Bitwise.scala 50:65:@3469.4]
  assign _T_4101 = _T_4070[30]; // @[Bitwise.scala 50:65:@3470.4]
  assign _T_4102 = _T_4070[31]; // @[Bitwise.scala 50:65:@3471.4]
  assign _T_4103 = _T_4071 + _T_4072; // @[Bitwise.scala 48:55:@3472.4]
  assign _T_4104 = _T_4073 + _T_4074; // @[Bitwise.scala 48:55:@3473.4]
  assign _T_4105 = _T_4103 + _T_4104; // @[Bitwise.scala 48:55:@3474.4]
  assign _T_4106 = _T_4075 + _T_4076; // @[Bitwise.scala 48:55:@3475.4]
  assign _T_4107 = _T_4077 + _T_4078; // @[Bitwise.scala 48:55:@3476.4]
  assign _T_4108 = _T_4106 + _T_4107; // @[Bitwise.scala 48:55:@3477.4]
  assign _T_4109 = _T_4105 + _T_4108; // @[Bitwise.scala 48:55:@3478.4]
  assign _T_4110 = _T_4079 + _T_4080; // @[Bitwise.scala 48:55:@3479.4]
  assign _T_4111 = _T_4081 + _T_4082; // @[Bitwise.scala 48:55:@3480.4]
  assign _T_4112 = _T_4110 + _T_4111; // @[Bitwise.scala 48:55:@3481.4]
  assign _T_4113 = _T_4083 + _T_4084; // @[Bitwise.scala 48:55:@3482.4]
  assign _T_4114 = _T_4085 + _T_4086; // @[Bitwise.scala 48:55:@3483.4]
  assign _T_4115 = _T_4113 + _T_4114; // @[Bitwise.scala 48:55:@3484.4]
  assign _T_4116 = _T_4112 + _T_4115; // @[Bitwise.scala 48:55:@3485.4]
  assign _T_4117 = _T_4109 + _T_4116; // @[Bitwise.scala 48:55:@3486.4]
  assign _T_4118 = _T_4087 + _T_4088; // @[Bitwise.scala 48:55:@3487.4]
  assign _T_4119 = _T_4089 + _T_4090; // @[Bitwise.scala 48:55:@3488.4]
  assign _T_4120 = _T_4118 + _T_4119; // @[Bitwise.scala 48:55:@3489.4]
  assign _T_4121 = _T_4091 + _T_4092; // @[Bitwise.scala 48:55:@3490.4]
  assign _T_4122 = _T_4093 + _T_4094; // @[Bitwise.scala 48:55:@3491.4]
  assign _T_4123 = _T_4121 + _T_4122; // @[Bitwise.scala 48:55:@3492.4]
  assign _T_4124 = _T_4120 + _T_4123; // @[Bitwise.scala 48:55:@3493.4]
  assign _T_4125 = _T_4095 + _T_4096; // @[Bitwise.scala 48:55:@3494.4]
  assign _T_4126 = _T_4097 + _T_4098; // @[Bitwise.scala 48:55:@3495.4]
  assign _T_4127 = _T_4125 + _T_4126; // @[Bitwise.scala 48:55:@3496.4]
  assign _T_4128 = _T_4099 + _T_4100; // @[Bitwise.scala 48:55:@3497.4]
  assign _T_4129 = _T_4101 + _T_4102; // @[Bitwise.scala 48:55:@3498.4]
  assign _T_4130 = _T_4128 + _T_4129; // @[Bitwise.scala 48:55:@3499.4]
  assign _T_4131 = _T_4127 + _T_4130; // @[Bitwise.scala 48:55:@3500.4]
  assign _T_4132 = _T_4124 + _T_4131; // @[Bitwise.scala 48:55:@3501.4]
  assign _T_4133 = _T_4117 + _T_4132; // @[Bitwise.scala 48:55:@3502.4]
  assign _T_4197 = _T_1124[32:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3567.4]
  assign _T_4198 = _T_4197[0]; // @[Bitwise.scala 50:65:@3568.4]
  assign _T_4199 = _T_4197[1]; // @[Bitwise.scala 50:65:@3569.4]
  assign _T_4200 = _T_4197[2]; // @[Bitwise.scala 50:65:@3570.4]
  assign _T_4201 = _T_4197[3]; // @[Bitwise.scala 50:65:@3571.4]
  assign _T_4202 = _T_4197[4]; // @[Bitwise.scala 50:65:@3572.4]
  assign _T_4203 = _T_4197[5]; // @[Bitwise.scala 50:65:@3573.4]
  assign _T_4204 = _T_4197[6]; // @[Bitwise.scala 50:65:@3574.4]
  assign _T_4205 = _T_4197[7]; // @[Bitwise.scala 50:65:@3575.4]
  assign _T_4206 = _T_4197[8]; // @[Bitwise.scala 50:65:@3576.4]
  assign _T_4207 = _T_4197[9]; // @[Bitwise.scala 50:65:@3577.4]
  assign _T_4208 = _T_4197[10]; // @[Bitwise.scala 50:65:@3578.4]
  assign _T_4209 = _T_4197[11]; // @[Bitwise.scala 50:65:@3579.4]
  assign _T_4210 = _T_4197[12]; // @[Bitwise.scala 50:65:@3580.4]
  assign _T_4211 = _T_4197[13]; // @[Bitwise.scala 50:65:@3581.4]
  assign _T_4212 = _T_4197[14]; // @[Bitwise.scala 50:65:@3582.4]
  assign _T_4213 = _T_4197[15]; // @[Bitwise.scala 50:65:@3583.4]
  assign _T_4214 = _T_4197[16]; // @[Bitwise.scala 50:65:@3584.4]
  assign _T_4215 = _T_4197[17]; // @[Bitwise.scala 50:65:@3585.4]
  assign _T_4216 = _T_4197[18]; // @[Bitwise.scala 50:65:@3586.4]
  assign _T_4217 = _T_4197[19]; // @[Bitwise.scala 50:65:@3587.4]
  assign _T_4218 = _T_4197[20]; // @[Bitwise.scala 50:65:@3588.4]
  assign _T_4219 = _T_4197[21]; // @[Bitwise.scala 50:65:@3589.4]
  assign _T_4220 = _T_4197[22]; // @[Bitwise.scala 50:65:@3590.4]
  assign _T_4221 = _T_4197[23]; // @[Bitwise.scala 50:65:@3591.4]
  assign _T_4222 = _T_4197[24]; // @[Bitwise.scala 50:65:@3592.4]
  assign _T_4223 = _T_4197[25]; // @[Bitwise.scala 50:65:@3593.4]
  assign _T_4224 = _T_4197[26]; // @[Bitwise.scala 50:65:@3594.4]
  assign _T_4225 = _T_4197[27]; // @[Bitwise.scala 50:65:@3595.4]
  assign _T_4226 = _T_4197[28]; // @[Bitwise.scala 50:65:@3596.4]
  assign _T_4227 = _T_4197[29]; // @[Bitwise.scala 50:65:@3597.4]
  assign _T_4228 = _T_4197[30]; // @[Bitwise.scala 50:65:@3598.4]
  assign _T_4229 = _T_4197[31]; // @[Bitwise.scala 50:65:@3599.4]
  assign _T_4230 = _T_4197[32]; // @[Bitwise.scala 50:65:@3600.4]
  assign _T_4231 = _T_4198 + _T_4199; // @[Bitwise.scala 48:55:@3601.4]
  assign _T_4232 = _T_4200 + _T_4201; // @[Bitwise.scala 48:55:@3602.4]
  assign _T_4233 = _T_4231 + _T_4232; // @[Bitwise.scala 48:55:@3603.4]
  assign _T_4234 = _T_4202 + _T_4203; // @[Bitwise.scala 48:55:@3604.4]
  assign _T_4235 = _T_4204 + _T_4205; // @[Bitwise.scala 48:55:@3605.4]
  assign _T_4236 = _T_4234 + _T_4235; // @[Bitwise.scala 48:55:@3606.4]
  assign _T_4237 = _T_4233 + _T_4236; // @[Bitwise.scala 48:55:@3607.4]
  assign _T_4238 = _T_4206 + _T_4207; // @[Bitwise.scala 48:55:@3608.4]
  assign _T_4239 = _T_4208 + _T_4209; // @[Bitwise.scala 48:55:@3609.4]
  assign _T_4240 = _T_4238 + _T_4239; // @[Bitwise.scala 48:55:@3610.4]
  assign _T_4241 = _T_4210 + _T_4211; // @[Bitwise.scala 48:55:@3611.4]
  assign _T_4242 = _T_4212 + _T_4213; // @[Bitwise.scala 48:55:@3612.4]
  assign _T_4243 = _T_4241 + _T_4242; // @[Bitwise.scala 48:55:@3613.4]
  assign _T_4244 = _T_4240 + _T_4243; // @[Bitwise.scala 48:55:@3614.4]
  assign _T_4245 = _T_4237 + _T_4244; // @[Bitwise.scala 48:55:@3615.4]
  assign _T_4246 = _T_4214 + _T_4215; // @[Bitwise.scala 48:55:@3616.4]
  assign _T_4247 = _T_4216 + _T_4217; // @[Bitwise.scala 48:55:@3617.4]
  assign _T_4248 = _T_4246 + _T_4247; // @[Bitwise.scala 48:55:@3618.4]
  assign _T_4249 = _T_4218 + _T_4219; // @[Bitwise.scala 48:55:@3619.4]
  assign _T_4250 = _T_4220 + _T_4221; // @[Bitwise.scala 48:55:@3620.4]
  assign _T_4251 = _T_4249 + _T_4250; // @[Bitwise.scala 48:55:@3621.4]
  assign _T_4252 = _T_4248 + _T_4251; // @[Bitwise.scala 48:55:@3622.4]
  assign _T_4253 = _T_4222 + _T_4223; // @[Bitwise.scala 48:55:@3623.4]
  assign _T_4254 = _T_4224 + _T_4225; // @[Bitwise.scala 48:55:@3624.4]
  assign _T_4255 = _T_4253 + _T_4254; // @[Bitwise.scala 48:55:@3625.4]
  assign _T_4256 = _T_4226 + _T_4227; // @[Bitwise.scala 48:55:@3626.4]
  assign _T_4257 = _T_4229 + _T_4230; // @[Bitwise.scala 48:55:@3627.4]
  assign _GEN_656 = {{1'd0}, _T_4228}; // @[Bitwise.scala 48:55:@3628.4]
  assign _T_4258 = _GEN_656 + _T_4257; // @[Bitwise.scala 48:55:@3628.4]
  assign _GEN_657 = {{1'd0}, _T_4256}; // @[Bitwise.scala 48:55:@3629.4]
  assign _T_4259 = _GEN_657 + _T_4258; // @[Bitwise.scala 48:55:@3629.4]
  assign _GEN_658 = {{1'd0}, _T_4255}; // @[Bitwise.scala 48:55:@3630.4]
  assign _T_4260 = _GEN_658 + _T_4259; // @[Bitwise.scala 48:55:@3630.4]
  assign _GEN_659 = {{1'd0}, _T_4252}; // @[Bitwise.scala 48:55:@3631.4]
  assign _T_4261 = _GEN_659 + _T_4260; // @[Bitwise.scala 48:55:@3631.4]
  assign _GEN_660 = {{1'd0}, _T_4245}; // @[Bitwise.scala 48:55:@3632.4]
  assign _T_4262 = _GEN_660 + _T_4261; // @[Bitwise.scala 48:55:@3632.4]
  assign _T_4326 = _T_1124[33:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3697.4]
  assign _T_4327 = _T_4326[0]; // @[Bitwise.scala 50:65:@3698.4]
  assign _T_4328 = _T_4326[1]; // @[Bitwise.scala 50:65:@3699.4]
  assign _T_4329 = _T_4326[2]; // @[Bitwise.scala 50:65:@3700.4]
  assign _T_4330 = _T_4326[3]; // @[Bitwise.scala 50:65:@3701.4]
  assign _T_4331 = _T_4326[4]; // @[Bitwise.scala 50:65:@3702.4]
  assign _T_4332 = _T_4326[5]; // @[Bitwise.scala 50:65:@3703.4]
  assign _T_4333 = _T_4326[6]; // @[Bitwise.scala 50:65:@3704.4]
  assign _T_4334 = _T_4326[7]; // @[Bitwise.scala 50:65:@3705.4]
  assign _T_4335 = _T_4326[8]; // @[Bitwise.scala 50:65:@3706.4]
  assign _T_4336 = _T_4326[9]; // @[Bitwise.scala 50:65:@3707.4]
  assign _T_4337 = _T_4326[10]; // @[Bitwise.scala 50:65:@3708.4]
  assign _T_4338 = _T_4326[11]; // @[Bitwise.scala 50:65:@3709.4]
  assign _T_4339 = _T_4326[12]; // @[Bitwise.scala 50:65:@3710.4]
  assign _T_4340 = _T_4326[13]; // @[Bitwise.scala 50:65:@3711.4]
  assign _T_4341 = _T_4326[14]; // @[Bitwise.scala 50:65:@3712.4]
  assign _T_4342 = _T_4326[15]; // @[Bitwise.scala 50:65:@3713.4]
  assign _T_4343 = _T_4326[16]; // @[Bitwise.scala 50:65:@3714.4]
  assign _T_4344 = _T_4326[17]; // @[Bitwise.scala 50:65:@3715.4]
  assign _T_4345 = _T_4326[18]; // @[Bitwise.scala 50:65:@3716.4]
  assign _T_4346 = _T_4326[19]; // @[Bitwise.scala 50:65:@3717.4]
  assign _T_4347 = _T_4326[20]; // @[Bitwise.scala 50:65:@3718.4]
  assign _T_4348 = _T_4326[21]; // @[Bitwise.scala 50:65:@3719.4]
  assign _T_4349 = _T_4326[22]; // @[Bitwise.scala 50:65:@3720.4]
  assign _T_4350 = _T_4326[23]; // @[Bitwise.scala 50:65:@3721.4]
  assign _T_4351 = _T_4326[24]; // @[Bitwise.scala 50:65:@3722.4]
  assign _T_4352 = _T_4326[25]; // @[Bitwise.scala 50:65:@3723.4]
  assign _T_4353 = _T_4326[26]; // @[Bitwise.scala 50:65:@3724.4]
  assign _T_4354 = _T_4326[27]; // @[Bitwise.scala 50:65:@3725.4]
  assign _T_4355 = _T_4326[28]; // @[Bitwise.scala 50:65:@3726.4]
  assign _T_4356 = _T_4326[29]; // @[Bitwise.scala 50:65:@3727.4]
  assign _T_4357 = _T_4326[30]; // @[Bitwise.scala 50:65:@3728.4]
  assign _T_4358 = _T_4326[31]; // @[Bitwise.scala 50:65:@3729.4]
  assign _T_4359 = _T_4326[32]; // @[Bitwise.scala 50:65:@3730.4]
  assign _T_4360 = _T_4326[33]; // @[Bitwise.scala 50:65:@3731.4]
  assign _T_4361 = _T_4327 + _T_4328; // @[Bitwise.scala 48:55:@3732.4]
  assign _T_4362 = _T_4329 + _T_4330; // @[Bitwise.scala 48:55:@3733.4]
  assign _T_4363 = _T_4361 + _T_4362; // @[Bitwise.scala 48:55:@3734.4]
  assign _T_4364 = _T_4331 + _T_4332; // @[Bitwise.scala 48:55:@3735.4]
  assign _T_4365 = _T_4333 + _T_4334; // @[Bitwise.scala 48:55:@3736.4]
  assign _T_4366 = _T_4364 + _T_4365; // @[Bitwise.scala 48:55:@3737.4]
  assign _T_4367 = _T_4363 + _T_4366; // @[Bitwise.scala 48:55:@3738.4]
  assign _T_4368 = _T_4335 + _T_4336; // @[Bitwise.scala 48:55:@3739.4]
  assign _T_4369 = _T_4337 + _T_4338; // @[Bitwise.scala 48:55:@3740.4]
  assign _T_4370 = _T_4368 + _T_4369; // @[Bitwise.scala 48:55:@3741.4]
  assign _T_4371 = _T_4339 + _T_4340; // @[Bitwise.scala 48:55:@3742.4]
  assign _T_4372 = _T_4342 + _T_4343; // @[Bitwise.scala 48:55:@3743.4]
  assign _GEN_661 = {{1'd0}, _T_4341}; // @[Bitwise.scala 48:55:@3744.4]
  assign _T_4373 = _GEN_661 + _T_4372; // @[Bitwise.scala 48:55:@3744.4]
  assign _GEN_662 = {{1'd0}, _T_4371}; // @[Bitwise.scala 48:55:@3745.4]
  assign _T_4374 = _GEN_662 + _T_4373; // @[Bitwise.scala 48:55:@3745.4]
  assign _GEN_663 = {{1'd0}, _T_4370}; // @[Bitwise.scala 48:55:@3746.4]
  assign _T_4375 = _GEN_663 + _T_4374; // @[Bitwise.scala 48:55:@3746.4]
  assign _GEN_664 = {{1'd0}, _T_4367}; // @[Bitwise.scala 48:55:@3747.4]
  assign _T_4376 = _GEN_664 + _T_4375; // @[Bitwise.scala 48:55:@3747.4]
  assign _T_4377 = _T_4344 + _T_4345; // @[Bitwise.scala 48:55:@3748.4]
  assign _T_4378 = _T_4346 + _T_4347; // @[Bitwise.scala 48:55:@3749.4]
  assign _T_4379 = _T_4377 + _T_4378; // @[Bitwise.scala 48:55:@3750.4]
  assign _T_4380 = _T_4348 + _T_4349; // @[Bitwise.scala 48:55:@3751.4]
  assign _T_4381 = _T_4350 + _T_4351; // @[Bitwise.scala 48:55:@3752.4]
  assign _T_4382 = _T_4380 + _T_4381; // @[Bitwise.scala 48:55:@3753.4]
  assign _T_4383 = _T_4379 + _T_4382; // @[Bitwise.scala 48:55:@3754.4]
  assign _T_4384 = _T_4352 + _T_4353; // @[Bitwise.scala 48:55:@3755.4]
  assign _T_4385 = _T_4354 + _T_4355; // @[Bitwise.scala 48:55:@3756.4]
  assign _T_4386 = _T_4384 + _T_4385; // @[Bitwise.scala 48:55:@3757.4]
  assign _T_4387 = _T_4356 + _T_4357; // @[Bitwise.scala 48:55:@3758.4]
  assign _T_4388 = _T_4359 + _T_4360; // @[Bitwise.scala 48:55:@3759.4]
  assign _GEN_665 = {{1'd0}, _T_4358}; // @[Bitwise.scala 48:55:@3760.4]
  assign _T_4389 = _GEN_665 + _T_4388; // @[Bitwise.scala 48:55:@3760.4]
  assign _GEN_666 = {{1'd0}, _T_4387}; // @[Bitwise.scala 48:55:@3761.4]
  assign _T_4390 = _GEN_666 + _T_4389; // @[Bitwise.scala 48:55:@3761.4]
  assign _GEN_667 = {{1'd0}, _T_4386}; // @[Bitwise.scala 48:55:@3762.4]
  assign _T_4391 = _GEN_667 + _T_4390; // @[Bitwise.scala 48:55:@3762.4]
  assign _GEN_668 = {{1'd0}, _T_4383}; // @[Bitwise.scala 48:55:@3763.4]
  assign _T_4392 = _GEN_668 + _T_4391; // @[Bitwise.scala 48:55:@3763.4]
  assign _T_4393 = _T_4376 + _T_4392; // @[Bitwise.scala 48:55:@3764.4]
  assign _T_4457 = _T_1124[34:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3829.4]
  assign _T_4458 = _T_4457[0]; // @[Bitwise.scala 50:65:@3830.4]
  assign _T_4459 = _T_4457[1]; // @[Bitwise.scala 50:65:@3831.4]
  assign _T_4460 = _T_4457[2]; // @[Bitwise.scala 50:65:@3832.4]
  assign _T_4461 = _T_4457[3]; // @[Bitwise.scala 50:65:@3833.4]
  assign _T_4462 = _T_4457[4]; // @[Bitwise.scala 50:65:@3834.4]
  assign _T_4463 = _T_4457[5]; // @[Bitwise.scala 50:65:@3835.4]
  assign _T_4464 = _T_4457[6]; // @[Bitwise.scala 50:65:@3836.4]
  assign _T_4465 = _T_4457[7]; // @[Bitwise.scala 50:65:@3837.4]
  assign _T_4466 = _T_4457[8]; // @[Bitwise.scala 50:65:@3838.4]
  assign _T_4467 = _T_4457[9]; // @[Bitwise.scala 50:65:@3839.4]
  assign _T_4468 = _T_4457[10]; // @[Bitwise.scala 50:65:@3840.4]
  assign _T_4469 = _T_4457[11]; // @[Bitwise.scala 50:65:@3841.4]
  assign _T_4470 = _T_4457[12]; // @[Bitwise.scala 50:65:@3842.4]
  assign _T_4471 = _T_4457[13]; // @[Bitwise.scala 50:65:@3843.4]
  assign _T_4472 = _T_4457[14]; // @[Bitwise.scala 50:65:@3844.4]
  assign _T_4473 = _T_4457[15]; // @[Bitwise.scala 50:65:@3845.4]
  assign _T_4474 = _T_4457[16]; // @[Bitwise.scala 50:65:@3846.4]
  assign _T_4475 = _T_4457[17]; // @[Bitwise.scala 50:65:@3847.4]
  assign _T_4476 = _T_4457[18]; // @[Bitwise.scala 50:65:@3848.4]
  assign _T_4477 = _T_4457[19]; // @[Bitwise.scala 50:65:@3849.4]
  assign _T_4478 = _T_4457[20]; // @[Bitwise.scala 50:65:@3850.4]
  assign _T_4479 = _T_4457[21]; // @[Bitwise.scala 50:65:@3851.4]
  assign _T_4480 = _T_4457[22]; // @[Bitwise.scala 50:65:@3852.4]
  assign _T_4481 = _T_4457[23]; // @[Bitwise.scala 50:65:@3853.4]
  assign _T_4482 = _T_4457[24]; // @[Bitwise.scala 50:65:@3854.4]
  assign _T_4483 = _T_4457[25]; // @[Bitwise.scala 50:65:@3855.4]
  assign _T_4484 = _T_4457[26]; // @[Bitwise.scala 50:65:@3856.4]
  assign _T_4485 = _T_4457[27]; // @[Bitwise.scala 50:65:@3857.4]
  assign _T_4486 = _T_4457[28]; // @[Bitwise.scala 50:65:@3858.4]
  assign _T_4487 = _T_4457[29]; // @[Bitwise.scala 50:65:@3859.4]
  assign _T_4488 = _T_4457[30]; // @[Bitwise.scala 50:65:@3860.4]
  assign _T_4489 = _T_4457[31]; // @[Bitwise.scala 50:65:@3861.4]
  assign _T_4490 = _T_4457[32]; // @[Bitwise.scala 50:65:@3862.4]
  assign _T_4491 = _T_4457[33]; // @[Bitwise.scala 50:65:@3863.4]
  assign _T_4492 = _T_4457[34]; // @[Bitwise.scala 50:65:@3864.4]
  assign _T_4493 = _T_4458 + _T_4459; // @[Bitwise.scala 48:55:@3865.4]
  assign _T_4494 = _T_4460 + _T_4461; // @[Bitwise.scala 48:55:@3866.4]
  assign _T_4495 = _T_4493 + _T_4494; // @[Bitwise.scala 48:55:@3867.4]
  assign _T_4496 = _T_4462 + _T_4463; // @[Bitwise.scala 48:55:@3868.4]
  assign _T_4497 = _T_4464 + _T_4465; // @[Bitwise.scala 48:55:@3869.4]
  assign _T_4498 = _T_4496 + _T_4497; // @[Bitwise.scala 48:55:@3870.4]
  assign _T_4499 = _T_4495 + _T_4498; // @[Bitwise.scala 48:55:@3871.4]
  assign _T_4500 = _T_4466 + _T_4467; // @[Bitwise.scala 48:55:@3872.4]
  assign _T_4501 = _T_4468 + _T_4469; // @[Bitwise.scala 48:55:@3873.4]
  assign _T_4502 = _T_4500 + _T_4501; // @[Bitwise.scala 48:55:@3874.4]
  assign _T_4503 = _T_4470 + _T_4471; // @[Bitwise.scala 48:55:@3875.4]
  assign _T_4504 = _T_4473 + _T_4474; // @[Bitwise.scala 48:55:@3876.4]
  assign _GEN_669 = {{1'd0}, _T_4472}; // @[Bitwise.scala 48:55:@3877.4]
  assign _T_4505 = _GEN_669 + _T_4504; // @[Bitwise.scala 48:55:@3877.4]
  assign _GEN_670 = {{1'd0}, _T_4503}; // @[Bitwise.scala 48:55:@3878.4]
  assign _T_4506 = _GEN_670 + _T_4505; // @[Bitwise.scala 48:55:@3878.4]
  assign _GEN_671 = {{1'd0}, _T_4502}; // @[Bitwise.scala 48:55:@3879.4]
  assign _T_4507 = _GEN_671 + _T_4506; // @[Bitwise.scala 48:55:@3879.4]
  assign _GEN_672 = {{1'd0}, _T_4499}; // @[Bitwise.scala 48:55:@3880.4]
  assign _T_4508 = _GEN_672 + _T_4507; // @[Bitwise.scala 48:55:@3880.4]
  assign _T_4509 = _T_4475 + _T_4476; // @[Bitwise.scala 48:55:@3881.4]
  assign _T_4510 = _T_4477 + _T_4478; // @[Bitwise.scala 48:55:@3882.4]
  assign _T_4511 = _T_4509 + _T_4510; // @[Bitwise.scala 48:55:@3883.4]
  assign _T_4512 = _T_4479 + _T_4480; // @[Bitwise.scala 48:55:@3884.4]
  assign _T_4513 = _T_4482 + _T_4483; // @[Bitwise.scala 48:55:@3885.4]
  assign _GEN_673 = {{1'd0}, _T_4481}; // @[Bitwise.scala 48:55:@3886.4]
  assign _T_4514 = _GEN_673 + _T_4513; // @[Bitwise.scala 48:55:@3886.4]
  assign _GEN_674 = {{1'd0}, _T_4512}; // @[Bitwise.scala 48:55:@3887.4]
  assign _T_4515 = _GEN_674 + _T_4514; // @[Bitwise.scala 48:55:@3887.4]
  assign _GEN_675 = {{1'd0}, _T_4511}; // @[Bitwise.scala 48:55:@3888.4]
  assign _T_4516 = _GEN_675 + _T_4515; // @[Bitwise.scala 48:55:@3888.4]
  assign _T_4517 = _T_4484 + _T_4485; // @[Bitwise.scala 48:55:@3889.4]
  assign _T_4518 = _T_4486 + _T_4487; // @[Bitwise.scala 48:55:@3890.4]
  assign _T_4519 = _T_4517 + _T_4518; // @[Bitwise.scala 48:55:@3891.4]
  assign _T_4520 = _T_4488 + _T_4489; // @[Bitwise.scala 48:55:@3892.4]
  assign _T_4521 = _T_4491 + _T_4492; // @[Bitwise.scala 48:55:@3893.4]
  assign _GEN_676 = {{1'd0}, _T_4490}; // @[Bitwise.scala 48:55:@3894.4]
  assign _T_4522 = _GEN_676 + _T_4521; // @[Bitwise.scala 48:55:@3894.4]
  assign _GEN_677 = {{1'd0}, _T_4520}; // @[Bitwise.scala 48:55:@3895.4]
  assign _T_4523 = _GEN_677 + _T_4522; // @[Bitwise.scala 48:55:@3895.4]
  assign _GEN_678 = {{1'd0}, _T_4519}; // @[Bitwise.scala 48:55:@3896.4]
  assign _T_4524 = _GEN_678 + _T_4523; // @[Bitwise.scala 48:55:@3896.4]
  assign _T_4525 = _T_4516 + _T_4524; // @[Bitwise.scala 48:55:@3897.4]
  assign _T_4526 = _T_4508 + _T_4525; // @[Bitwise.scala 48:55:@3898.4]
  assign _T_4590 = _T_1124[35:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@3963.4]
  assign _T_4591 = _T_4590[0]; // @[Bitwise.scala 50:65:@3964.4]
  assign _T_4592 = _T_4590[1]; // @[Bitwise.scala 50:65:@3965.4]
  assign _T_4593 = _T_4590[2]; // @[Bitwise.scala 50:65:@3966.4]
  assign _T_4594 = _T_4590[3]; // @[Bitwise.scala 50:65:@3967.4]
  assign _T_4595 = _T_4590[4]; // @[Bitwise.scala 50:65:@3968.4]
  assign _T_4596 = _T_4590[5]; // @[Bitwise.scala 50:65:@3969.4]
  assign _T_4597 = _T_4590[6]; // @[Bitwise.scala 50:65:@3970.4]
  assign _T_4598 = _T_4590[7]; // @[Bitwise.scala 50:65:@3971.4]
  assign _T_4599 = _T_4590[8]; // @[Bitwise.scala 50:65:@3972.4]
  assign _T_4600 = _T_4590[9]; // @[Bitwise.scala 50:65:@3973.4]
  assign _T_4601 = _T_4590[10]; // @[Bitwise.scala 50:65:@3974.4]
  assign _T_4602 = _T_4590[11]; // @[Bitwise.scala 50:65:@3975.4]
  assign _T_4603 = _T_4590[12]; // @[Bitwise.scala 50:65:@3976.4]
  assign _T_4604 = _T_4590[13]; // @[Bitwise.scala 50:65:@3977.4]
  assign _T_4605 = _T_4590[14]; // @[Bitwise.scala 50:65:@3978.4]
  assign _T_4606 = _T_4590[15]; // @[Bitwise.scala 50:65:@3979.4]
  assign _T_4607 = _T_4590[16]; // @[Bitwise.scala 50:65:@3980.4]
  assign _T_4608 = _T_4590[17]; // @[Bitwise.scala 50:65:@3981.4]
  assign _T_4609 = _T_4590[18]; // @[Bitwise.scala 50:65:@3982.4]
  assign _T_4610 = _T_4590[19]; // @[Bitwise.scala 50:65:@3983.4]
  assign _T_4611 = _T_4590[20]; // @[Bitwise.scala 50:65:@3984.4]
  assign _T_4612 = _T_4590[21]; // @[Bitwise.scala 50:65:@3985.4]
  assign _T_4613 = _T_4590[22]; // @[Bitwise.scala 50:65:@3986.4]
  assign _T_4614 = _T_4590[23]; // @[Bitwise.scala 50:65:@3987.4]
  assign _T_4615 = _T_4590[24]; // @[Bitwise.scala 50:65:@3988.4]
  assign _T_4616 = _T_4590[25]; // @[Bitwise.scala 50:65:@3989.4]
  assign _T_4617 = _T_4590[26]; // @[Bitwise.scala 50:65:@3990.4]
  assign _T_4618 = _T_4590[27]; // @[Bitwise.scala 50:65:@3991.4]
  assign _T_4619 = _T_4590[28]; // @[Bitwise.scala 50:65:@3992.4]
  assign _T_4620 = _T_4590[29]; // @[Bitwise.scala 50:65:@3993.4]
  assign _T_4621 = _T_4590[30]; // @[Bitwise.scala 50:65:@3994.4]
  assign _T_4622 = _T_4590[31]; // @[Bitwise.scala 50:65:@3995.4]
  assign _T_4623 = _T_4590[32]; // @[Bitwise.scala 50:65:@3996.4]
  assign _T_4624 = _T_4590[33]; // @[Bitwise.scala 50:65:@3997.4]
  assign _T_4625 = _T_4590[34]; // @[Bitwise.scala 50:65:@3998.4]
  assign _T_4626 = _T_4590[35]; // @[Bitwise.scala 50:65:@3999.4]
  assign _T_4627 = _T_4591 + _T_4592; // @[Bitwise.scala 48:55:@4000.4]
  assign _T_4628 = _T_4593 + _T_4594; // @[Bitwise.scala 48:55:@4001.4]
  assign _T_4629 = _T_4627 + _T_4628; // @[Bitwise.scala 48:55:@4002.4]
  assign _T_4630 = _T_4595 + _T_4596; // @[Bitwise.scala 48:55:@4003.4]
  assign _T_4631 = _T_4598 + _T_4599; // @[Bitwise.scala 48:55:@4004.4]
  assign _GEN_679 = {{1'd0}, _T_4597}; // @[Bitwise.scala 48:55:@4005.4]
  assign _T_4632 = _GEN_679 + _T_4631; // @[Bitwise.scala 48:55:@4005.4]
  assign _GEN_680 = {{1'd0}, _T_4630}; // @[Bitwise.scala 48:55:@4006.4]
  assign _T_4633 = _GEN_680 + _T_4632; // @[Bitwise.scala 48:55:@4006.4]
  assign _GEN_681 = {{1'd0}, _T_4629}; // @[Bitwise.scala 48:55:@4007.4]
  assign _T_4634 = _GEN_681 + _T_4633; // @[Bitwise.scala 48:55:@4007.4]
  assign _T_4635 = _T_4600 + _T_4601; // @[Bitwise.scala 48:55:@4008.4]
  assign _T_4636 = _T_4602 + _T_4603; // @[Bitwise.scala 48:55:@4009.4]
  assign _T_4637 = _T_4635 + _T_4636; // @[Bitwise.scala 48:55:@4010.4]
  assign _T_4638 = _T_4604 + _T_4605; // @[Bitwise.scala 48:55:@4011.4]
  assign _T_4639 = _T_4607 + _T_4608; // @[Bitwise.scala 48:55:@4012.4]
  assign _GEN_682 = {{1'd0}, _T_4606}; // @[Bitwise.scala 48:55:@4013.4]
  assign _T_4640 = _GEN_682 + _T_4639; // @[Bitwise.scala 48:55:@4013.4]
  assign _GEN_683 = {{1'd0}, _T_4638}; // @[Bitwise.scala 48:55:@4014.4]
  assign _T_4641 = _GEN_683 + _T_4640; // @[Bitwise.scala 48:55:@4014.4]
  assign _GEN_684 = {{1'd0}, _T_4637}; // @[Bitwise.scala 48:55:@4015.4]
  assign _T_4642 = _GEN_684 + _T_4641; // @[Bitwise.scala 48:55:@4015.4]
  assign _T_4643 = _T_4634 + _T_4642; // @[Bitwise.scala 48:55:@4016.4]
  assign _T_4644 = _T_4609 + _T_4610; // @[Bitwise.scala 48:55:@4017.4]
  assign _T_4645 = _T_4611 + _T_4612; // @[Bitwise.scala 48:55:@4018.4]
  assign _T_4646 = _T_4644 + _T_4645; // @[Bitwise.scala 48:55:@4019.4]
  assign _T_4647 = _T_4613 + _T_4614; // @[Bitwise.scala 48:55:@4020.4]
  assign _T_4648 = _T_4616 + _T_4617; // @[Bitwise.scala 48:55:@4021.4]
  assign _GEN_685 = {{1'd0}, _T_4615}; // @[Bitwise.scala 48:55:@4022.4]
  assign _T_4649 = _GEN_685 + _T_4648; // @[Bitwise.scala 48:55:@4022.4]
  assign _GEN_686 = {{1'd0}, _T_4647}; // @[Bitwise.scala 48:55:@4023.4]
  assign _T_4650 = _GEN_686 + _T_4649; // @[Bitwise.scala 48:55:@4023.4]
  assign _GEN_687 = {{1'd0}, _T_4646}; // @[Bitwise.scala 48:55:@4024.4]
  assign _T_4651 = _GEN_687 + _T_4650; // @[Bitwise.scala 48:55:@4024.4]
  assign _T_4652 = _T_4618 + _T_4619; // @[Bitwise.scala 48:55:@4025.4]
  assign _T_4653 = _T_4620 + _T_4621; // @[Bitwise.scala 48:55:@4026.4]
  assign _T_4654 = _T_4652 + _T_4653; // @[Bitwise.scala 48:55:@4027.4]
  assign _T_4655 = _T_4622 + _T_4623; // @[Bitwise.scala 48:55:@4028.4]
  assign _T_4656 = _T_4625 + _T_4626; // @[Bitwise.scala 48:55:@4029.4]
  assign _GEN_688 = {{1'd0}, _T_4624}; // @[Bitwise.scala 48:55:@4030.4]
  assign _T_4657 = _GEN_688 + _T_4656; // @[Bitwise.scala 48:55:@4030.4]
  assign _GEN_689 = {{1'd0}, _T_4655}; // @[Bitwise.scala 48:55:@4031.4]
  assign _T_4658 = _GEN_689 + _T_4657; // @[Bitwise.scala 48:55:@4031.4]
  assign _GEN_690 = {{1'd0}, _T_4654}; // @[Bitwise.scala 48:55:@4032.4]
  assign _T_4659 = _GEN_690 + _T_4658; // @[Bitwise.scala 48:55:@4032.4]
  assign _T_4660 = _T_4651 + _T_4659; // @[Bitwise.scala 48:55:@4033.4]
  assign _T_4661 = _T_4643 + _T_4660; // @[Bitwise.scala 48:55:@4034.4]
  assign _T_4725 = _T_1124[36:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4099.4]
  assign _T_4726 = _T_4725[0]; // @[Bitwise.scala 50:65:@4100.4]
  assign _T_4727 = _T_4725[1]; // @[Bitwise.scala 50:65:@4101.4]
  assign _T_4728 = _T_4725[2]; // @[Bitwise.scala 50:65:@4102.4]
  assign _T_4729 = _T_4725[3]; // @[Bitwise.scala 50:65:@4103.4]
  assign _T_4730 = _T_4725[4]; // @[Bitwise.scala 50:65:@4104.4]
  assign _T_4731 = _T_4725[5]; // @[Bitwise.scala 50:65:@4105.4]
  assign _T_4732 = _T_4725[6]; // @[Bitwise.scala 50:65:@4106.4]
  assign _T_4733 = _T_4725[7]; // @[Bitwise.scala 50:65:@4107.4]
  assign _T_4734 = _T_4725[8]; // @[Bitwise.scala 50:65:@4108.4]
  assign _T_4735 = _T_4725[9]; // @[Bitwise.scala 50:65:@4109.4]
  assign _T_4736 = _T_4725[10]; // @[Bitwise.scala 50:65:@4110.4]
  assign _T_4737 = _T_4725[11]; // @[Bitwise.scala 50:65:@4111.4]
  assign _T_4738 = _T_4725[12]; // @[Bitwise.scala 50:65:@4112.4]
  assign _T_4739 = _T_4725[13]; // @[Bitwise.scala 50:65:@4113.4]
  assign _T_4740 = _T_4725[14]; // @[Bitwise.scala 50:65:@4114.4]
  assign _T_4741 = _T_4725[15]; // @[Bitwise.scala 50:65:@4115.4]
  assign _T_4742 = _T_4725[16]; // @[Bitwise.scala 50:65:@4116.4]
  assign _T_4743 = _T_4725[17]; // @[Bitwise.scala 50:65:@4117.4]
  assign _T_4744 = _T_4725[18]; // @[Bitwise.scala 50:65:@4118.4]
  assign _T_4745 = _T_4725[19]; // @[Bitwise.scala 50:65:@4119.4]
  assign _T_4746 = _T_4725[20]; // @[Bitwise.scala 50:65:@4120.4]
  assign _T_4747 = _T_4725[21]; // @[Bitwise.scala 50:65:@4121.4]
  assign _T_4748 = _T_4725[22]; // @[Bitwise.scala 50:65:@4122.4]
  assign _T_4749 = _T_4725[23]; // @[Bitwise.scala 50:65:@4123.4]
  assign _T_4750 = _T_4725[24]; // @[Bitwise.scala 50:65:@4124.4]
  assign _T_4751 = _T_4725[25]; // @[Bitwise.scala 50:65:@4125.4]
  assign _T_4752 = _T_4725[26]; // @[Bitwise.scala 50:65:@4126.4]
  assign _T_4753 = _T_4725[27]; // @[Bitwise.scala 50:65:@4127.4]
  assign _T_4754 = _T_4725[28]; // @[Bitwise.scala 50:65:@4128.4]
  assign _T_4755 = _T_4725[29]; // @[Bitwise.scala 50:65:@4129.4]
  assign _T_4756 = _T_4725[30]; // @[Bitwise.scala 50:65:@4130.4]
  assign _T_4757 = _T_4725[31]; // @[Bitwise.scala 50:65:@4131.4]
  assign _T_4758 = _T_4725[32]; // @[Bitwise.scala 50:65:@4132.4]
  assign _T_4759 = _T_4725[33]; // @[Bitwise.scala 50:65:@4133.4]
  assign _T_4760 = _T_4725[34]; // @[Bitwise.scala 50:65:@4134.4]
  assign _T_4761 = _T_4725[35]; // @[Bitwise.scala 50:65:@4135.4]
  assign _T_4762 = _T_4725[36]; // @[Bitwise.scala 50:65:@4136.4]
  assign _T_4763 = _T_4726 + _T_4727; // @[Bitwise.scala 48:55:@4137.4]
  assign _T_4764 = _T_4728 + _T_4729; // @[Bitwise.scala 48:55:@4138.4]
  assign _T_4765 = _T_4763 + _T_4764; // @[Bitwise.scala 48:55:@4139.4]
  assign _T_4766 = _T_4730 + _T_4731; // @[Bitwise.scala 48:55:@4140.4]
  assign _T_4767 = _T_4733 + _T_4734; // @[Bitwise.scala 48:55:@4141.4]
  assign _GEN_691 = {{1'd0}, _T_4732}; // @[Bitwise.scala 48:55:@4142.4]
  assign _T_4768 = _GEN_691 + _T_4767; // @[Bitwise.scala 48:55:@4142.4]
  assign _GEN_692 = {{1'd0}, _T_4766}; // @[Bitwise.scala 48:55:@4143.4]
  assign _T_4769 = _GEN_692 + _T_4768; // @[Bitwise.scala 48:55:@4143.4]
  assign _GEN_693 = {{1'd0}, _T_4765}; // @[Bitwise.scala 48:55:@4144.4]
  assign _T_4770 = _GEN_693 + _T_4769; // @[Bitwise.scala 48:55:@4144.4]
  assign _T_4771 = _T_4735 + _T_4736; // @[Bitwise.scala 48:55:@4145.4]
  assign _T_4772 = _T_4737 + _T_4738; // @[Bitwise.scala 48:55:@4146.4]
  assign _T_4773 = _T_4771 + _T_4772; // @[Bitwise.scala 48:55:@4147.4]
  assign _T_4774 = _T_4739 + _T_4740; // @[Bitwise.scala 48:55:@4148.4]
  assign _T_4775 = _T_4742 + _T_4743; // @[Bitwise.scala 48:55:@4149.4]
  assign _GEN_694 = {{1'd0}, _T_4741}; // @[Bitwise.scala 48:55:@4150.4]
  assign _T_4776 = _GEN_694 + _T_4775; // @[Bitwise.scala 48:55:@4150.4]
  assign _GEN_695 = {{1'd0}, _T_4774}; // @[Bitwise.scala 48:55:@4151.4]
  assign _T_4777 = _GEN_695 + _T_4776; // @[Bitwise.scala 48:55:@4151.4]
  assign _GEN_696 = {{1'd0}, _T_4773}; // @[Bitwise.scala 48:55:@4152.4]
  assign _T_4778 = _GEN_696 + _T_4777; // @[Bitwise.scala 48:55:@4152.4]
  assign _T_4779 = _T_4770 + _T_4778; // @[Bitwise.scala 48:55:@4153.4]
  assign _T_4780 = _T_4744 + _T_4745; // @[Bitwise.scala 48:55:@4154.4]
  assign _T_4781 = _T_4746 + _T_4747; // @[Bitwise.scala 48:55:@4155.4]
  assign _T_4782 = _T_4780 + _T_4781; // @[Bitwise.scala 48:55:@4156.4]
  assign _T_4783 = _T_4748 + _T_4749; // @[Bitwise.scala 48:55:@4157.4]
  assign _T_4784 = _T_4751 + _T_4752; // @[Bitwise.scala 48:55:@4158.4]
  assign _GEN_697 = {{1'd0}, _T_4750}; // @[Bitwise.scala 48:55:@4159.4]
  assign _T_4785 = _GEN_697 + _T_4784; // @[Bitwise.scala 48:55:@4159.4]
  assign _GEN_698 = {{1'd0}, _T_4783}; // @[Bitwise.scala 48:55:@4160.4]
  assign _T_4786 = _GEN_698 + _T_4785; // @[Bitwise.scala 48:55:@4160.4]
  assign _GEN_699 = {{1'd0}, _T_4782}; // @[Bitwise.scala 48:55:@4161.4]
  assign _T_4787 = _GEN_699 + _T_4786; // @[Bitwise.scala 48:55:@4161.4]
  assign _T_4788 = _T_4753 + _T_4754; // @[Bitwise.scala 48:55:@4162.4]
  assign _T_4789 = _T_4756 + _T_4757; // @[Bitwise.scala 48:55:@4163.4]
  assign _GEN_700 = {{1'd0}, _T_4755}; // @[Bitwise.scala 48:55:@4164.4]
  assign _T_4790 = _GEN_700 + _T_4789; // @[Bitwise.scala 48:55:@4164.4]
  assign _GEN_701 = {{1'd0}, _T_4788}; // @[Bitwise.scala 48:55:@4165.4]
  assign _T_4791 = _GEN_701 + _T_4790; // @[Bitwise.scala 48:55:@4165.4]
  assign _T_4792 = _T_4758 + _T_4759; // @[Bitwise.scala 48:55:@4166.4]
  assign _T_4793 = _T_4761 + _T_4762; // @[Bitwise.scala 48:55:@4167.4]
  assign _GEN_702 = {{1'd0}, _T_4760}; // @[Bitwise.scala 48:55:@4168.4]
  assign _T_4794 = _GEN_702 + _T_4793; // @[Bitwise.scala 48:55:@4168.4]
  assign _GEN_703 = {{1'd0}, _T_4792}; // @[Bitwise.scala 48:55:@4169.4]
  assign _T_4795 = _GEN_703 + _T_4794; // @[Bitwise.scala 48:55:@4169.4]
  assign _T_4796 = _T_4791 + _T_4795; // @[Bitwise.scala 48:55:@4170.4]
  assign _T_4797 = _T_4787 + _T_4796; // @[Bitwise.scala 48:55:@4171.4]
  assign _T_4798 = _T_4779 + _T_4797; // @[Bitwise.scala 48:55:@4172.4]
  assign _T_4862 = _T_1124[37:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4237.4]
  assign _T_4863 = _T_4862[0]; // @[Bitwise.scala 50:65:@4238.4]
  assign _T_4864 = _T_4862[1]; // @[Bitwise.scala 50:65:@4239.4]
  assign _T_4865 = _T_4862[2]; // @[Bitwise.scala 50:65:@4240.4]
  assign _T_4866 = _T_4862[3]; // @[Bitwise.scala 50:65:@4241.4]
  assign _T_4867 = _T_4862[4]; // @[Bitwise.scala 50:65:@4242.4]
  assign _T_4868 = _T_4862[5]; // @[Bitwise.scala 50:65:@4243.4]
  assign _T_4869 = _T_4862[6]; // @[Bitwise.scala 50:65:@4244.4]
  assign _T_4870 = _T_4862[7]; // @[Bitwise.scala 50:65:@4245.4]
  assign _T_4871 = _T_4862[8]; // @[Bitwise.scala 50:65:@4246.4]
  assign _T_4872 = _T_4862[9]; // @[Bitwise.scala 50:65:@4247.4]
  assign _T_4873 = _T_4862[10]; // @[Bitwise.scala 50:65:@4248.4]
  assign _T_4874 = _T_4862[11]; // @[Bitwise.scala 50:65:@4249.4]
  assign _T_4875 = _T_4862[12]; // @[Bitwise.scala 50:65:@4250.4]
  assign _T_4876 = _T_4862[13]; // @[Bitwise.scala 50:65:@4251.4]
  assign _T_4877 = _T_4862[14]; // @[Bitwise.scala 50:65:@4252.4]
  assign _T_4878 = _T_4862[15]; // @[Bitwise.scala 50:65:@4253.4]
  assign _T_4879 = _T_4862[16]; // @[Bitwise.scala 50:65:@4254.4]
  assign _T_4880 = _T_4862[17]; // @[Bitwise.scala 50:65:@4255.4]
  assign _T_4881 = _T_4862[18]; // @[Bitwise.scala 50:65:@4256.4]
  assign _T_4882 = _T_4862[19]; // @[Bitwise.scala 50:65:@4257.4]
  assign _T_4883 = _T_4862[20]; // @[Bitwise.scala 50:65:@4258.4]
  assign _T_4884 = _T_4862[21]; // @[Bitwise.scala 50:65:@4259.4]
  assign _T_4885 = _T_4862[22]; // @[Bitwise.scala 50:65:@4260.4]
  assign _T_4886 = _T_4862[23]; // @[Bitwise.scala 50:65:@4261.4]
  assign _T_4887 = _T_4862[24]; // @[Bitwise.scala 50:65:@4262.4]
  assign _T_4888 = _T_4862[25]; // @[Bitwise.scala 50:65:@4263.4]
  assign _T_4889 = _T_4862[26]; // @[Bitwise.scala 50:65:@4264.4]
  assign _T_4890 = _T_4862[27]; // @[Bitwise.scala 50:65:@4265.4]
  assign _T_4891 = _T_4862[28]; // @[Bitwise.scala 50:65:@4266.4]
  assign _T_4892 = _T_4862[29]; // @[Bitwise.scala 50:65:@4267.4]
  assign _T_4893 = _T_4862[30]; // @[Bitwise.scala 50:65:@4268.4]
  assign _T_4894 = _T_4862[31]; // @[Bitwise.scala 50:65:@4269.4]
  assign _T_4895 = _T_4862[32]; // @[Bitwise.scala 50:65:@4270.4]
  assign _T_4896 = _T_4862[33]; // @[Bitwise.scala 50:65:@4271.4]
  assign _T_4897 = _T_4862[34]; // @[Bitwise.scala 50:65:@4272.4]
  assign _T_4898 = _T_4862[35]; // @[Bitwise.scala 50:65:@4273.4]
  assign _T_4899 = _T_4862[36]; // @[Bitwise.scala 50:65:@4274.4]
  assign _T_4900 = _T_4862[37]; // @[Bitwise.scala 50:65:@4275.4]
  assign _T_4901 = _T_4863 + _T_4864; // @[Bitwise.scala 48:55:@4276.4]
  assign _T_4902 = _T_4865 + _T_4866; // @[Bitwise.scala 48:55:@4277.4]
  assign _T_4903 = _T_4901 + _T_4902; // @[Bitwise.scala 48:55:@4278.4]
  assign _T_4904 = _T_4867 + _T_4868; // @[Bitwise.scala 48:55:@4279.4]
  assign _T_4905 = _T_4870 + _T_4871; // @[Bitwise.scala 48:55:@4280.4]
  assign _GEN_704 = {{1'd0}, _T_4869}; // @[Bitwise.scala 48:55:@4281.4]
  assign _T_4906 = _GEN_704 + _T_4905; // @[Bitwise.scala 48:55:@4281.4]
  assign _GEN_705 = {{1'd0}, _T_4904}; // @[Bitwise.scala 48:55:@4282.4]
  assign _T_4907 = _GEN_705 + _T_4906; // @[Bitwise.scala 48:55:@4282.4]
  assign _GEN_706 = {{1'd0}, _T_4903}; // @[Bitwise.scala 48:55:@4283.4]
  assign _T_4908 = _GEN_706 + _T_4907; // @[Bitwise.scala 48:55:@4283.4]
  assign _T_4909 = _T_4872 + _T_4873; // @[Bitwise.scala 48:55:@4284.4]
  assign _T_4910 = _T_4875 + _T_4876; // @[Bitwise.scala 48:55:@4285.4]
  assign _GEN_707 = {{1'd0}, _T_4874}; // @[Bitwise.scala 48:55:@4286.4]
  assign _T_4911 = _GEN_707 + _T_4910; // @[Bitwise.scala 48:55:@4286.4]
  assign _GEN_708 = {{1'd0}, _T_4909}; // @[Bitwise.scala 48:55:@4287.4]
  assign _T_4912 = _GEN_708 + _T_4911; // @[Bitwise.scala 48:55:@4287.4]
  assign _T_4913 = _T_4877 + _T_4878; // @[Bitwise.scala 48:55:@4288.4]
  assign _T_4914 = _T_4880 + _T_4881; // @[Bitwise.scala 48:55:@4289.4]
  assign _GEN_709 = {{1'd0}, _T_4879}; // @[Bitwise.scala 48:55:@4290.4]
  assign _T_4915 = _GEN_709 + _T_4914; // @[Bitwise.scala 48:55:@4290.4]
  assign _GEN_710 = {{1'd0}, _T_4913}; // @[Bitwise.scala 48:55:@4291.4]
  assign _T_4916 = _GEN_710 + _T_4915; // @[Bitwise.scala 48:55:@4291.4]
  assign _T_4917 = _T_4912 + _T_4916; // @[Bitwise.scala 48:55:@4292.4]
  assign _T_4918 = _T_4908 + _T_4917; // @[Bitwise.scala 48:55:@4293.4]
  assign _T_4919 = _T_4882 + _T_4883; // @[Bitwise.scala 48:55:@4294.4]
  assign _T_4920 = _T_4884 + _T_4885; // @[Bitwise.scala 48:55:@4295.4]
  assign _T_4921 = _T_4919 + _T_4920; // @[Bitwise.scala 48:55:@4296.4]
  assign _T_4922 = _T_4886 + _T_4887; // @[Bitwise.scala 48:55:@4297.4]
  assign _T_4923 = _T_4889 + _T_4890; // @[Bitwise.scala 48:55:@4298.4]
  assign _GEN_711 = {{1'd0}, _T_4888}; // @[Bitwise.scala 48:55:@4299.4]
  assign _T_4924 = _GEN_711 + _T_4923; // @[Bitwise.scala 48:55:@4299.4]
  assign _GEN_712 = {{1'd0}, _T_4922}; // @[Bitwise.scala 48:55:@4300.4]
  assign _T_4925 = _GEN_712 + _T_4924; // @[Bitwise.scala 48:55:@4300.4]
  assign _GEN_713 = {{1'd0}, _T_4921}; // @[Bitwise.scala 48:55:@4301.4]
  assign _T_4926 = _GEN_713 + _T_4925; // @[Bitwise.scala 48:55:@4301.4]
  assign _T_4927 = _T_4891 + _T_4892; // @[Bitwise.scala 48:55:@4302.4]
  assign _T_4928 = _T_4894 + _T_4895; // @[Bitwise.scala 48:55:@4303.4]
  assign _GEN_714 = {{1'd0}, _T_4893}; // @[Bitwise.scala 48:55:@4304.4]
  assign _T_4929 = _GEN_714 + _T_4928; // @[Bitwise.scala 48:55:@4304.4]
  assign _GEN_715 = {{1'd0}, _T_4927}; // @[Bitwise.scala 48:55:@4305.4]
  assign _T_4930 = _GEN_715 + _T_4929; // @[Bitwise.scala 48:55:@4305.4]
  assign _T_4931 = _T_4896 + _T_4897; // @[Bitwise.scala 48:55:@4306.4]
  assign _T_4932 = _T_4899 + _T_4900; // @[Bitwise.scala 48:55:@4307.4]
  assign _GEN_716 = {{1'd0}, _T_4898}; // @[Bitwise.scala 48:55:@4308.4]
  assign _T_4933 = _GEN_716 + _T_4932; // @[Bitwise.scala 48:55:@4308.4]
  assign _GEN_717 = {{1'd0}, _T_4931}; // @[Bitwise.scala 48:55:@4309.4]
  assign _T_4934 = _GEN_717 + _T_4933; // @[Bitwise.scala 48:55:@4309.4]
  assign _T_4935 = _T_4930 + _T_4934; // @[Bitwise.scala 48:55:@4310.4]
  assign _T_4936 = _T_4926 + _T_4935; // @[Bitwise.scala 48:55:@4311.4]
  assign _T_4937 = _T_4918 + _T_4936; // @[Bitwise.scala 48:55:@4312.4]
  assign _T_5001 = _T_1124[38:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4377.4]
  assign _T_5002 = _T_5001[0]; // @[Bitwise.scala 50:65:@4378.4]
  assign _T_5003 = _T_5001[1]; // @[Bitwise.scala 50:65:@4379.4]
  assign _T_5004 = _T_5001[2]; // @[Bitwise.scala 50:65:@4380.4]
  assign _T_5005 = _T_5001[3]; // @[Bitwise.scala 50:65:@4381.4]
  assign _T_5006 = _T_5001[4]; // @[Bitwise.scala 50:65:@4382.4]
  assign _T_5007 = _T_5001[5]; // @[Bitwise.scala 50:65:@4383.4]
  assign _T_5008 = _T_5001[6]; // @[Bitwise.scala 50:65:@4384.4]
  assign _T_5009 = _T_5001[7]; // @[Bitwise.scala 50:65:@4385.4]
  assign _T_5010 = _T_5001[8]; // @[Bitwise.scala 50:65:@4386.4]
  assign _T_5011 = _T_5001[9]; // @[Bitwise.scala 50:65:@4387.4]
  assign _T_5012 = _T_5001[10]; // @[Bitwise.scala 50:65:@4388.4]
  assign _T_5013 = _T_5001[11]; // @[Bitwise.scala 50:65:@4389.4]
  assign _T_5014 = _T_5001[12]; // @[Bitwise.scala 50:65:@4390.4]
  assign _T_5015 = _T_5001[13]; // @[Bitwise.scala 50:65:@4391.4]
  assign _T_5016 = _T_5001[14]; // @[Bitwise.scala 50:65:@4392.4]
  assign _T_5017 = _T_5001[15]; // @[Bitwise.scala 50:65:@4393.4]
  assign _T_5018 = _T_5001[16]; // @[Bitwise.scala 50:65:@4394.4]
  assign _T_5019 = _T_5001[17]; // @[Bitwise.scala 50:65:@4395.4]
  assign _T_5020 = _T_5001[18]; // @[Bitwise.scala 50:65:@4396.4]
  assign _T_5021 = _T_5001[19]; // @[Bitwise.scala 50:65:@4397.4]
  assign _T_5022 = _T_5001[20]; // @[Bitwise.scala 50:65:@4398.4]
  assign _T_5023 = _T_5001[21]; // @[Bitwise.scala 50:65:@4399.4]
  assign _T_5024 = _T_5001[22]; // @[Bitwise.scala 50:65:@4400.4]
  assign _T_5025 = _T_5001[23]; // @[Bitwise.scala 50:65:@4401.4]
  assign _T_5026 = _T_5001[24]; // @[Bitwise.scala 50:65:@4402.4]
  assign _T_5027 = _T_5001[25]; // @[Bitwise.scala 50:65:@4403.4]
  assign _T_5028 = _T_5001[26]; // @[Bitwise.scala 50:65:@4404.4]
  assign _T_5029 = _T_5001[27]; // @[Bitwise.scala 50:65:@4405.4]
  assign _T_5030 = _T_5001[28]; // @[Bitwise.scala 50:65:@4406.4]
  assign _T_5031 = _T_5001[29]; // @[Bitwise.scala 50:65:@4407.4]
  assign _T_5032 = _T_5001[30]; // @[Bitwise.scala 50:65:@4408.4]
  assign _T_5033 = _T_5001[31]; // @[Bitwise.scala 50:65:@4409.4]
  assign _T_5034 = _T_5001[32]; // @[Bitwise.scala 50:65:@4410.4]
  assign _T_5035 = _T_5001[33]; // @[Bitwise.scala 50:65:@4411.4]
  assign _T_5036 = _T_5001[34]; // @[Bitwise.scala 50:65:@4412.4]
  assign _T_5037 = _T_5001[35]; // @[Bitwise.scala 50:65:@4413.4]
  assign _T_5038 = _T_5001[36]; // @[Bitwise.scala 50:65:@4414.4]
  assign _T_5039 = _T_5001[37]; // @[Bitwise.scala 50:65:@4415.4]
  assign _T_5040 = _T_5001[38]; // @[Bitwise.scala 50:65:@4416.4]
  assign _T_5041 = _T_5002 + _T_5003; // @[Bitwise.scala 48:55:@4417.4]
  assign _T_5042 = _T_5004 + _T_5005; // @[Bitwise.scala 48:55:@4418.4]
  assign _T_5043 = _T_5041 + _T_5042; // @[Bitwise.scala 48:55:@4419.4]
  assign _T_5044 = _T_5006 + _T_5007; // @[Bitwise.scala 48:55:@4420.4]
  assign _T_5045 = _T_5009 + _T_5010; // @[Bitwise.scala 48:55:@4421.4]
  assign _GEN_718 = {{1'd0}, _T_5008}; // @[Bitwise.scala 48:55:@4422.4]
  assign _T_5046 = _GEN_718 + _T_5045; // @[Bitwise.scala 48:55:@4422.4]
  assign _GEN_719 = {{1'd0}, _T_5044}; // @[Bitwise.scala 48:55:@4423.4]
  assign _T_5047 = _GEN_719 + _T_5046; // @[Bitwise.scala 48:55:@4423.4]
  assign _GEN_720 = {{1'd0}, _T_5043}; // @[Bitwise.scala 48:55:@4424.4]
  assign _T_5048 = _GEN_720 + _T_5047; // @[Bitwise.scala 48:55:@4424.4]
  assign _T_5049 = _T_5011 + _T_5012; // @[Bitwise.scala 48:55:@4425.4]
  assign _T_5050 = _T_5014 + _T_5015; // @[Bitwise.scala 48:55:@4426.4]
  assign _GEN_721 = {{1'd0}, _T_5013}; // @[Bitwise.scala 48:55:@4427.4]
  assign _T_5051 = _GEN_721 + _T_5050; // @[Bitwise.scala 48:55:@4427.4]
  assign _GEN_722 = {{1'd0}, _T_5049}; // @[Bitwise.scala 48:55:@4428.4]
  assign _T_5052 = _GEN_722 + _T_5051; // @[Bitwise.scala 48:55:@4428.4]
  assign _T_5053 = _T_5016 + _T_5017; // @[Bitwise.scala 48:55:@4429.4]
  assign _T_5054 = _T_5019 + _T_5020; // @[Bitwise.scala 48:55:@4430.4]
  assign _GEN_723 = {{1'd0}, _T_5018}; // @[Bitwise.scala 48:55:@4431.4]
  assign _T_5055 = _GEN_723 + _T_5054; // @[Bitwise.scala 48:55:@4431.4]
  assign _GEN_724 = {{1'd0}, _T_5053}; // @[Bitwise.scala 48:55:@4432.4]
  assign _T_5056 = _GEN_724 + _T_5055; // @[Bitwise.scala 48:55:@4432.4]
  assign _T_5057 = _T_5052 + _T_5056; // @[Bitwise.scala 48:55:@4433.4]
  assign _T_5058 = _T_5048 + _T_5057; // @[Bitwise.scala 48:55:@4434.4]
  assign _T_5059 = _T_5021 + _T_5022; // @[Bitwise.scala 48:55:@4435.4]
  assign _T_5060 = _T_5024 + _T_5025; // @[Bitwise.scala 48:55:@4436.4]
  assign _GEN_725 = {{1'd0}, _T_5023}; // @[Bitwise.scala 48:55:@4437.4]
  assign _T_5061 = _GEN_725 + _T_5060; // @[Bitwise.scala 48:55:@4437.4]
  assign _GEN_726 = {{1'd0}, _T_5059}; // @[Bitwise.scala 48:55:@4438.4]
  assign _T_5062 = _GEN_726 + _T_5061; // @[Bitwise.scala 48:55:@4438.4]
  assign _T_5063 = _T_5026 + _T_5027; // @[Bitwise.scala 48:55:@4439.4]
  assign _T_5064 = _T_5029 + _T_5030; // @[Bitwise.scala 48:55:@4440.4]
  assign _GEN_727 = {{1'd0}, _T_5028}; // @[Bitwise.scala 48:55:@4441.4]
  assign _T_5065 = _GEN_727 + _T_5064; // @[Bitwise.scala 48:55:@4441.4]
  assign _GEN_728 = {{1'd0}, _T_5063}; // @[Bitwise.scala 48:55:@4442.4]
  assign _T_5066 = _GEN_728 + _T_5065; // @[Bitwise.scala 48:55:@4442.4]
  assign _T_5067 = _T_5062 + _T_5066; // @[Bitwise.scala 48:55:@4443.4]
  assign _T_5068 = _T_5031 + _T_5032; // @[Bitwise.scala 48:55:@4444.4]
  assign _T_5069 = _T_5034 + _T_5035; // @[Bitwise.scala 48:55:@4445.4]
  assign _GEN_729 = {{1'd0}, _T_5033}; // @[Bitwise.scala 48:55:@4446.4]
  assign _T_5070 = _GEN_729 + _T_5069; // @[Bitwise.scala 48:55:@4446.4]
  assign _GEN_730 = {{1'd0}, _T_5068}; // @[Bitwise.scala 48:55:@4447.4]
  assign _T_5071 = _GEN_730 + _T_5070; // @[Bitwise.scala 48:55:@4447.4]
  assign _T_5072 = _T_5036 + _T_5037; // @[Bitwise.scala 48:55:@4448.4]
  assign _T_5073 = _T_5039 + _T_5040; // @[Bitwise.scala 48:55:@4449.4]
  assign _GEN_731 = {{1'd0}, _T_5038}; // @[Bitwise.scala 48:55:@4450.4]
  assign _T_5074 = _GEN_731 + _T_5073; // @[Bitwise.scala 48:55:@4450.4]
  assign _GEN_732 = {{1'd0}, _T_5072}; // @[Bitwise.scala 48:55:@4451.4]
  assign _T_5075 = _GEN_732 + _T_5074; // @[Bitwise.scala 48:55:@4451.4]
  assign _T_5076 = _T_5071 + _T_5075; // @[Bitwise.scala 48:55:@4452.4]
  assign _T_5077 = _T_5067 + _T_5076; // @[Bitwise.scala 48:55:@4453.4]
  assign _T_5078 = _T_5058 + _T_5077; // @[Bitwise.scala 48:55:@4454.4]
  assign _T_5142 = _T_1124[39:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4519.4]
  assign _T_5143 = _T_5142[0]; // @[Bitwise.scala 50:65:@4520.4]
  assign _T_5144 = _T_5142[1]; // @[Bitwise.scala 50:65:@4521.4]
  assign _T_5145 = _T_5142[2]; // @[Bitwise.scala 50:65:@4522.4]
  assign _T_5146 = _T_5142[3]; // @[Bitwise.scala 50:65:@4523.4]
  assign _T_5147 = _T_5142[4]; // @[Bitwise.scala 50:65:@4524.4]
  assign _T_5148 = _T_5142[5]; // @[Bitwise.scala 50:65:@4525.4]
  assign _T_5149 = _T_5142[6]; // @[Bitwise.scala 50:65:@4526.4]
  assign _T_5150 = _T_5142[7]; // @[Bitwise.scala 50:65:@4527.4]
  assign _T_5151 = _T_5142[8]; // @[Bitwise.scala 50:65:@4528.4]
  assign _T_5152 = _T_5142[9]; // @[Bitwise.scala 50:65:@4529.4]
  assign _T_5153 = _T_5142[10]; // @[Bitwise.scala 50:65:@4530.4]
  assign _T_5154 = _T_5142[11]; // @[Bitwise.scala 50:65:@4531.4]
  assign _T_5155 = _T_5142[12]; // @[Bitwise.scala 50:65:@4532.4]
  assign _T_5156 = _T_5142[13]; // @[Bitwise.scala 50:65:@4533.4]
  assign _T_5157 = _T_5142[14]; // @[Bitwise.scala 50:65:@4534.4]
  assign _T_5158 = _T_5142[15]; // @[Bitwise.scala 50:65:@4535.4]
  assign _T_5159 = _T_5142[16]; // @[Bitwise.scala 50:65:@4536.4]
  assign _T_5160 = _T_5142[17]; // @[Bitwise.scala 50:65:@4537.4]
  assign _T_5161 = _T_5142[18]; // @[Bitwise.scala 50:65:@4538.4]
  assign _T_5162 = _T_5142[19]; // @[Bitwise.scala 50:65:@4539.4]
  assign _T_5163 = _T_5142[20]; // @[Bitwise.scala 50:65:@4540.4]
  assign _T_5164 = _T_5142[21]; // @[Bitwise.scala 50:65:@4541.4]
  assign _T_5165 = _T_5142[22]; // @[Bitwise.scala 50:65:@4542.4]
  assign _T_5166 = _T_5142[23]; // @[Bitwise.scala 50:65:@4543.4]
  assign _T_5167 = _T_5142[24]; // @[Bitwise.scala 50:65:@4544.4]
  assign _T_5168 = _T_5142[25]; // @[Bitwise.scala 50:65:@4545.4]
  assign _T_5169 = _T_5142[26]; // @[Bitwise.scala 50:65:@4546.4]
  assign _T_5170 = _T_5142[27]; // @[Bitwise.scala 50:65:@4547.4]
  assign _T_5171 = _T_5142[28]; // @[Bitwise.scala 50:65:@4548.4]
  assign _T_5172 = _T_5142[29]; // @[Bitwise.scala 50:65:@4549.4]
  assign _T_5173 = _T_5142[30]; // @[Bitwise.scala 50:65:@4550.4]
  assign _T_5174 = _T_5142[31]; // @[Bitwise.scala 50:65:@4551.4]
  assign _T_5175 = _T_5142[32]; // @[Bitwise.scala 50:65:@4552.4]
  assign _T_5176 = _T_5142[33]; // @[Bitwise.scala 50:65:@4553.4]
  assign _T_5177 = _T_5142[34]; // @[Bitwise.scala 50:65:@4554.4]
  assign _T_5178 = _T_5142[35]; // @[Bitwise.scala 50:65:@4555.4]
  assign _T_5179 = _T_5142[36]; // @[Bitwise.scala 50:65:@4556.4]
  assign _T_5180 = _T_5142[37]; // @[Bitwise.scala 50:65:@4557.4]
  assign _T_5181 = _T_5142[38]; // @[Bitwise.scala 50:65:@4558.4]
  assign _T_5182 = _T_5142[39]; // @[Bitwise.scala 50:65:@4559.4]
  assign _T_5183 = _T_5143 + _T_5144; // @[Bitwise.scala 48:55:@4560.4]
  assign _T_5184 = _T_5146 + _T_5147; // @[Bitwise.scala 48:55:@4561.4]
  assign _GEN_733 = {{1'd0}, _T_5145}; // @[Bitwise.scala 48:55:@4562.4]
  assign _T_5185 = _GEN_733 + _T_5184; // @[Bitwise.scala 48:55:@4562.4]
  assign _GEN_734 = {{1'd0}, _T_5183}; // @[Bitwise.scala 48:55:@4563.4]
  assign _T_5186 = _GEN_734 + _T_5185; // @[Bitwise.scala 48:55:@4563.4]
  assign _T_5187 = _T_5148 + _T_5149; // @[Bitwise.scala 48:55:@4564.4]
  assign _T_5188 = _T_5151 + _T_5152; // @[Bitwise.scala 48:55:@4565.4]
  assign _GEN_735 = {{1'd0}, _T_5150}; // @[Bitwise.scala 48:55:@4566.4]
  assign _T_5189 = _GEN_735 + _T_5188; // @[Bitwise.scala 48:55:@4566.4]
  assign _GEN_736 = {{1'd0}, _T_5187}; // @[Bitwise.scala 48:55:@4567.4]
  assign _T_5190 = _GEN_736 + _T_5189; // @[Bitwise.scala 48:55:@4567.4]
  assign _T_5191 = _T_5186 + _T_5190; // @[Bitwise.scala 48:55:@4568.4]
  assign _T_5192 = _T_5153 + _T_5154; // @[Bitwise.scala 48:55:@4569.4]
  assign _T_5193 = _T_5156 + _T_5157; // @[Bitwise.scala 48:55:@4570.4]
  assign _GEN_737 = {{1'd0}, _T_5155}; // @[Bitwise.scala 48:55:@4571.4]
  assign _T_5194 = _GEN_737 + _T_5193; // @[Bitwise.scala 48:55:@4571.4]
  assign _GEN_738 = {{1'd0}, _T_5192}; // @[Bitwise.scala 48:55:@4572.4]
  assign _T_5195 = _GEN_738 + _T_5194; // @[Bitwise.scala 48:55:@4572.4]
  assign _T_5196 = _T_5158 + _T_5159; // @[Bitwise.scala 48:55:@4573.4]
  assign _T_5197 = _T_5161 + _T_5162; // @[Bitwise.scala 48:55:@4574.4]
  assign _GEN_739 = {{1'd0}, _T_5160}; // @[Bitwise.scala 48:55:@4575.4]
  assign _T_5198 = _GEN_739 + _T_5197; // @[Bitwise.scala 48:55:@4575.4]
  assign _GEN_740 = {{1'd0}, _T_5196}; // @[Bitwise.scala 48:55:@4576.4]
  assign _T_5199 = _GEN_740 + _T_5198; // @[Bitwise.scala 48:55:@4576.4]
  assign _T_5200 = _T_5195 + _T_5199; // @[Bitwise.scala 48:55:@4577.4]
  assign _T_5201 = _T_5191 + _T_5200; // @[Bitwise.scala 48:55:@4578.4]
  assign _T_5202 = _T_5163 + _T_5164; // @[Bitwise.scala 48:55:@4579.4]
  assign _T_5203 = _T_5166 + _T_5167; // @[Bitwise.scala 48:55:@4580.4]
  assign _GEN_741 = {{1'd0}, _T_5165}; // @[Bitwise.scala 48:55:@4581.4]
  assign _T_5204 = _GEN_741 + _T_5203; // @[Bitwise.scala 48:55:@4581.4]
  assign _GEN_742 = {{1'd0}, _T_5202}; // @[Bitwise.scala 48:55:@4582.4]
  assign _T_5205 = _GEN_742 + _T_5204; // @[Bitwise.scala 48:55:@4582.4]
  assign _T_5206 = _T_5168 + _T_5169; // @[Bitwise.scala 48:55:@4583.4]
  assign _T_5207 = _T_5171 + _T_5172; // @[Bitwise.scala 48:55:@4584.4]
  assign _GEN_743 = {{1'd0}, _T_5170}; // @[Bitwise.scala 48:55:@4585.4]
  assign _T_5208 = _GEN_743 + _T_5207; // @[Bitwise.scala 48:55:@4585.4]
  assign _GEN_744 = {{1'd0}, _T_5206}; // @[Bitwise.scala 48:55:@4586.4]
  assign _T_5209 = _GEN_744 + _T_5208; // @[Bitwise.scala 48:55:@4586.4]
  assign _T_5210 = _T_5205 + _T_5209; // @[Bitwise.scala 48:55:@4587.4]
  assign _T_5211 = _T_5173 + _T_5174; // @[Bitwise.scala 48:55:@4588.4]
  assign _T_5212 = _T_5176 + _T_5177; // @[Bitwise.scala 48:55:@4589.4]
  assign _GEN_745 = {{1'd0}, _T_5175}; // @[Bitwise.scala 48:55:@4590.4]
  assign _T_5213 = _GEN_745 + _T_5212; // @[Bitwise.scala 48:55:@4590.4]
  assign _GEN_746 = {{1'd0}, _T_5211}; // @[Bitwise.scala 48:55:@4591.4]
  assign _T_5214 = _GEN_746 + _T_5213; // @[Bitwise.scala 48:55:@4591.4]
  assign _T_5215 = _T_5178 + _T_5179; // @[Bitwise.scala 48:55:@4592.4]
  assign _T_5216 = _T_5181 + _T_5182; // @[Bitwise.scala 48:55:@4593.4]
  assign _GEN_747 = {{1'd0}, _T_5180}; // @[Bitwise.scala 48:55:@4594.4]
  assign _T_5217 = _GEN_747 + _T_5216; // @[Bitwise.scala 48:55:@4594.4]
  assign _GEN_748 = {{1'd0}, _T_5215}; // @[Bitwise.scala 48:55:@4595.4]
  assign _T_5218 = _GEN_748 + _T_5217; // @[Bitwise.scala 48:55:@4595.4]
  assign _T_5219 = _T_5214 + _T_5218; // @[Bitwise.scala 48:55:@4596.4]
  assign _T_5220 = _T_5210 + _T_5219; // @[Bitwise.scala 48:55:@4597.4]
  assign _T_5221 = _T_5201 + _T_5220; // @[Bitwise.scala 48:55:@4598.4]
  assign _T_5285 = _T_1124[40:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4663.4]
  assign _T_5286 = _T_5285[0]; // @[Bitwise.scala 50:65:@4664.4]
  assign _T_5287 = _T_5285[1]; // @[Bitwise.scala 50:65:@4665.4]
  assign _T_5288 = _T_5285[2]; // @[Bitwise.scala 50:65:@4666.4]
  assign _T_5289 = _T_5285[3]; // @[Bitwise.scala 50:65:@4667.4]
  assign _T_5290 = _T_5285[4]; // @[Bitwise.scala 50:65:@4668.4]
  assign _T_5291 = _T_5285[5]; // @[Bitwise.scala 50:65:@4669.4]
  assign _T_5292 = _T_5285[6]; // @[Bitwise.scala 50:65:@4670.4]
  assign _T_5293 = _T_5285[7]; // @[Bitwise.scala 50:65:@4671.4]
  assign _T_5294 = _T_5285[8]; // @[Bitwise.scala 50:65:@4672.4]
  assign _T_5295 = _T_5285[9]; // @[Bitwise.scala 50:65:@4673.4]
  assign _T_5296 = _T_5285[10]; // @[Bitwise.scala 50:65:@4674.4]
  assign _T_5297 = _T_5285[11]; // @[Bitwise.scala 50:65:@4675.4]
  assign _T_5298 = _T_5285[12]; // @[Bitwise.scala 50:65:@4676.4]
  assign _T_5299 = _T_5285[13]; // @[Bitwise.scala 50:65:@4677.4]
  assign _T_5300 = _T_5285[14]; // @[Bitwise.scala 50:65:@4678.4]
  assign _T_5301 = _T_5285[15]; // @[Bitwise.scala 50:65:@4679.4]
  assign _T_5302 = _T_5285[16]; // @[Bitwise.scala 50:65:@4680.4]
  assign _T_5303 = _T_5285[17]; // @[Bitwise.scala 50:65:@4681.4]
  assign _T_5304 = _T_5285[18]; // @[Bitwise.scala 50:65:@4682.4]
  assign _T_5305 = _T_5285[19]; // @[Bitwise.scala 50:65:@4683.4]
  assign _T_5306 = _T_5285[20]; // @[Bitwise.scala 50:65:@4684.4]
  assign _T_5307 = _T_5285[21]; // @[Bitwise.scala 50:65:@4685.4]
  assign _T_5308 = _T_5285[22]; // @[Bitwise.scala 50:65:@4686.4]
  assign _T_5309 = _T_5285[23]; // @[Bitwise.scala 50:65:@4687.4]
  assign _T_5310 = _T_5285[24]; // @[Bitwise.scala 50:65:@4688.4]
  assign _T_5311 = _T_5285[25]; // @[Bitwise.scala 50:65:@4689.4]
  assign _T_5312 = _T_5285[26]; // @[Bitwise.scala 50:65:@4690.4]
  assign _T_5313 = _T_5285[27]; // @[Bitwise.scala 50:65:@4691.4]
  assign _T_5314 = _T_5285[28]; // @[Bitwise.scala 50:65:@4692.4]
  assign _T_5315 = _T_5285[29]; // @[Bitwise.scala 50:65:@4693.4]
  assign _T_5316 = _T_5285[30]; // @[Bitwise.scala 50:65:@4694.4]
  assign _T_5317 = _T_5285[31]; // @[Bitwise.scala 50:65:@4695.4]
  assign _T_5318 = _T_5285[32]; // @[Bitwise.scala 50:65:@4696.4]
  assign _T_5319 = _T_5285[33]; // @[Bitwise.scala 50:65:@4697.4]
  assign _T_5320 = _T_5285[34]; // @[Bitwise.scala 50:65:@4698.4]
  assign _T_5321 = _T_5285[35]; // @[Bitwise.scala 50:65:@4699.4]
  assign _T_5322 = _T_5285[36]; // @[Bitwise.scala 50:65:@4700.4]
  assign _T_5323 = _T_5285[37]; // @[Bitwise.scala 50:65:@4701.4]
  assign _T_5324 = _T_5285[38]; // @[Bitwise.scala 50:65:@4702.4]
  assign _T_5325 = _T_5285[39]; // @[Bitwise.scala 50:65:@4703.4]
  assign _T_5326 = _T_5285[40]; // @[Bitwise.scala 50:65:@4704.4]
  assign _T_5327 = _T_5286 + _T_5287; // @[Bitwise.scala 48:55:@4705.4]
  assign _T_5328 = _T_5289 + _T_5290; // @[Bitwise.scala 48:55:@4706.4]
  assign _GEN_749 = {{1'd0}, _T_5288}; // @[Bitwise.scala 48:55:@4707.4]
  assign _T_5329 = _GEN_749 + _T_5328; // @[Bitwise.scala 48:55:@4707.4]
  assign _GEN_750 = {{1'd0}, _T_5327}; // @[Bitwise.scala 48:55:@4708.4]
  assign _T_5330 = _GEN_750 + _T_5329; // @[Bitwise.scala 48:55:@4708.4]
  assign _T_5331 = _T_5291 + _T_5292; // @[Bitwise.scala 48:55:@4709.4]
  assign _T_5332 = _T_5294 + _T_5295; // @[Bitwise.scala 48:55:@4710.4]
  assign _GEN_751 = {{1'd0}, _T_5293}; // @[Bitwise.scala 48:55:@4711.4]
  assign _T_5333 = _GEN_751 + _T_5332; // @[Bitwise.scala 48:55:@4711.4]
  assign _GEN_752 = {{1'd0}, _T_5331}; // @[Bitwise.scala 48:55:@4712.4]
  assign _T_5334 = _GEN_752 + _T_5333; // @[Bitwise.scala 48:55:@4712.4]
  assign _T_5335 = _T_5330 + _T_5334; // @[Bitwise.scala 48:55:@4713.4]
  assign _T_5336 = _T_5296 + _T_5297; // @[Bitwise.scala 48:55:@4714.4]
  assign _T_5337 = _T_5299 + _T_5300; // @[Bitwise.scala 48:55:@4715.4]
  assign _GEN_753 = {{1'd0}, _T_5298}; // @[Bitwise.scala 48:55:@4716.4]
  assign _T_5338 = _GEN_753 + _T_5337; // @[Bitwise.scala 48:55:@4716.4]
  assign _GEN_754 = {{1'd0}, _T_5336}; // @[Bitwise.scala 48:55:@4717.4]
  assign _T_5339 = _GEN_754 + _T_5338; // @[Bitwise.scala 48:55:@4717.4]
  assign _T_5340 = _T_5301 + _T_5302; // @[Bitwise.scala 48:55:@4718.4]
  assign _T_5341 = _T_5304 + _T_5305; // @[Bitwise.scala 48:55:@4719.4]
  assign _GEN_755 = {{1'd0}, _T_5303}; // @[Bitwise.scala 48:55:@4720.4]
  assign _T_5342 = _GEN_755 + _T_5341; // @[Bitwise.scala 48:55:@4720.4]
  assign _GEN_756 = {{1'd0}, _T_5340}; // @[Bitwise.scala 48:55:@4721.4]
  assign _T_5343 = _GEN_756 + _T_5342; // @[Bitwise.scala 48:55:@4721.4]
  assign _T_5344 = _T_5339 + _T_5343; // @[Bitwise.scala 48:55:@4722.4]
  assign _T_5345 = _T_5335 + _T_5344; // @[Bitwise.scala 48:55:@4723.4]
  assign _T_5346 = _T_5306 + _T_5307; // @[Bitwise.scala 48:55:@4724.4]
  assign _T_5347 = _T_5309 + _T_5310; // @[Bitwise.scala 48:55:@4725.4]
  assign _GEN_757 = {{1'd0}, _T_5308}; // @[Bitwise.scala 48:55:@4726.4]
  assign _T_5348 = _GEN_757 + _T_5347; // @[Bitwise.scala 48:55:@4726.4]
  assign _GEN_758 = {{1'd0}, _T_5346}; // @[Bitwise.scala 48:55:@4727.4]
  assign _T_5349 = _GEN_758 + _T_5348; // @[Bitwise.scala 48:55:@4727.4]
  assign _T_5350 = _T_5311 + _T_5312; // @[Bitwise.scala 48:55:@4728.4]
  assign _T_5351 = _T_5314 + _T_5315; // @[Bitwise.scala 48:55:@4729.4]
  assign _GEN_759 = {{1'd0}, _T_5313}; // @[Bitwise.scala 48:55:@4730.4]
  assign _T_5352 = _GEN_759 + _T_5351; // @[Bitwise.scala 48:55:@4730.4]
  assign _GEN_760 = {{1'd0}, _T_5350}; // @[Bitwise.scala 48:55:@4731.4]
  assign _T_5353 = _GEN_760 + _T_5352; // @[Bitwise.scala 48:55:@4731.4]
  assign _T_5354 = _T_5349 + _T_5353; // @[Bitwise.scala 48:55:@4732.4]
  assign _T_5355 = _T_5316 + _T_5317; // @[Bitwise.scala 48:55:@4733.4]
  assign _T_5356 = _T_5319 + _T_5320; // @[Bitwise.scala 48:55:@4734.4]
  assign _GEN_761 = {{1'd0}, _T_5318}; // @[Bitwise.scala 48:55:@4735.4]
  assign _T_5357 = _GEN_761 + _T_5356; // @[Bitwise.scala 48:55:@4735.4]
  assign _GEN_762 = {{1'd0}, _T_5355}; // @[Bitwise.scala 48:55:@4736.4]
  assign _T_5358 = _GEN_762 + _T_5357; // @[Bitwise.scala 48:55:@4736.4]
  assign _T_5359 = _T_5322 + _T_5323; // @[Bitwise.scala 48:55:@4737.4]
  assign _GEN_763 = {{1'd0}, _T_5321}; // @[Bitwise.scala 48:55:@4738.4]
  assign _T_5360 = _GEN_763 + _T_5359; // @[Bitwise.scala 48:55:@4738.4]
  assign _T_5361 = _T_5325 + _T_5326; // @[Bitwise.scala 48:55:@4739.4]
  assign _GEN_764 = {{1'd0}, _T_5324}; // @[Bitwise.scala 48:55:@4740.4]
  assign _T_5362 = _GEN_764 + _T_5361; // @[Bitwise.scala 48:55:@4740.4]
  assign _T_5363 = _T_5360 + _T_5362; // @[Bitwise.scala 48:55:@4741.4]
  assign _T_5364 = _T_5358 + _T_5363; // @[Bitwise.scala 48:55:@4742.4]
  assign _T_5365 = _T_5354 + _T_5364; // @[Bitwise.scala 48:55:@4743.4]
  assign _T_5366 = _T_5345 + _T_5365; // @[Bitwise.scala 48:55:@4744.4]
  assign _T_5430 = _T_1124[41:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4809.4]
  assign _T_5431 = _T_5430[0]; // @[Bitwise.scala 50:65:@4810.4]
  assign _T_5432 = _T_5430[1]; // @[Bitwise.scala 50:65:@4811.4]
  assign _T_5433 = _T_5430[2]; // @[Bitwise.scala 50:65:@4812.4]
  assign _T_5434 = _T_5430[3]; // @[Bitwise.scala 50:65:@4813.4]
  assign _T_5435 = _T_5430[4]; // @[Bitwise.scala 50:65:@4814.4]
  assign _T_5436 = _T_5430[5]; // @[Bitwise.scala 50:65:@4815.4]
  assign _T_5437 = _T_5430[6]; // @[Bitwise.scala 50:65:@4816.4]
  assign _T_5438 = _T_5430[7]; // @[Bitwise.scala 50:65:@4817.4]
  assign _T_5439 = _T_5430[8]; // @[Bitwise.scala 50:65:@4818.4]
  assign _T_5440 = _T_5430[9]; // @[Bitwise.scala 50:65:@4819.4]
  assign _T_5441 = _T_5430[10]; // @[Bitwise.scala 50:65:@4820.4]
  assign _T_5442 = _T_5430[11]; // @[Bitwise.scala 50:65:@4821.4]
  assign _T_5443 = _T_5430[12]; // @[Bitwise.scala 50:65:@4822.4]
  assign _T_5444 = _T_5430[13]; // @[Bitwise.scala 50:65:@4823.4]
  assign _T_5445 = _T_5430[14]; // @[Bitwise.scala 50:65:@4824.4]
  assign _T_5446 = _T_5430[15]; // @[Bitwise.scala 50:65:@4825.4]
  assign _T_5447 = _T_5430[16]; // @[Bitwise.scala 50:65:@4826.4]
  assign _T_5448 = _T_5430[17]; // @[Bitwise.scala 50:65:@4827.4]
  assign _T_5449 = _T_5430[18]; // @[Bitwise.scala 50:65:@4828.4]
  assign _T_5450 = _T_5430[19]; // @[Bitwise.scala 50:65:@4829.4]
  assign _T_5451 = _T_5430[20]; // @[Bitwise.scala 50:65:@4830.4]
  assign _T_5452 = _T_5430[21]; // @[Bitwise.scala 50:65:@4831.4]
  assign _T_5453 = _T_5430[22]; // @[Bitwise.scala 50:65:@4832.4]
  assign _T_5454 = _T_5430[23]; // @[Bitwise.scala 50:65:@4833.4]
  assign _T_5455 = _T_5430[24]; // @[Bitwise.scala 50:65:@4834.4]
  assign _T_5456 = _T_5430[25]; // @[Bitwise.scala 50:65:@4835.4]
  assign _T_5457 = _T_5430[26]; // @[Bitwise.scala 50:65:@4836.4]
  assign _T_5458 = _T_5430[27]; // @[Bitwise.scala 50:65:@4837.4]
  assign _T_5459 = _T_5430[28]; // @[Bitwise.scala 50:65:@4838.4]
  assign _T_5460 = _T_5430[29]; // @[Bitwise.scala 50:65:@4839.4]
  assign _T_5461 = _T_5430[30]; // @[Bitwise.scala 50:65:@4840.4]
  assign _T_5462 = _T_5430[31]; // @[Bitwise.scala 50:65:@4841.4]
  assign _T_5463 = _T_5430[32]; // @[Bitwise.scala 50:65:@4842.4]
  assign _T_5464 = _T_5430[33]; // @[Bitwise.scala 50:65:@4843.4]
  assign _T_5465 = _T_5430[34]; // @[Bitwise.scala 50:65:@4844.4]
  assign _T_5466 = _T_5430[35]; // @[Bitwise.scala 50:65:@4845.4]
  assign _T_5467 = _T_5430[36]; // @[Bitwise.scala 50:65:@4846.4]
  assign _T_5468 = _T_5430[37]; // @[Bitwise.scala 50:65:@4847.4]
  assign _T_5469 = _T_5430[38]; // @[Bitwise.scala 50:65:@4848.4]
  assign _T_5470 = _T_5430[39]; // @[Bitwise.scala 50:65:@4849.4]
  assign _T_5471 = _T_5430[40]; // @[Bitwise.scala 50:65:@4850.4]
  assign _T_5472 = _T_5430[41]; // @[Bitwise.scala 50:65:@4851.4]
  assign _T_5473 = _T_5431 + _T_5432; // @[Bitwise.scala 48:55:@4852.4]
  assign _T_5474 = _T_5434 + _T_5435; // @[Bitwise.scala 48:55:@4853.4]
  assign _GEN_765 = {{1'd0}, _T_5433}; // @[Bitwise.scala 48:55:@4854.4]
  assign _T_5475 = _GEN_765 + _T_5474; // @[Bitwise.scala 48:55:@4854.4]
  assign _GEN_766 = {{1'd0}, _T_5473}; // @[Bitwise.scala 48:55:@4855.4]
  assign _T_5476 = _GEN_766 + _T_5475; // @[Bitwise.scala 48:55:@4855.4]
  assign _T_5477 = _T_5436 + _T_5437; // @[Bitwise.scala 48:55:@4856.4]
  assign _T_5478 = _T_5439 + _T_5440; // @[Bitwise.scala 48:55:@4857.4]
  assign _GEN_767 = {{1'd0}, _T_5438}; // @[Bitwise.scala 48:55:@4858.4]
  assign _T_5479 = _GEN_767 + _T_5478; // @[Bitwise.scala 48:55:@4858.4]
  assign _GEN_768 = {{1'd0}, _T_5477}; // @[Bitwise.scala 48:55:@4859.4]
  assign _T_5480 = _GEN_768 + _T_5479; // @[Bitwise.scala 48:55:@4859.4]
  assign _T_5481 = _T_5476 + _T_5480; // @[Bitwise.scala 48:55:@4860.4]
  assign _T_5482 = _T_5441 + _T_5442; // @[Bitwise.scala 48:55:@4861.4]
  assign _T_5483 = _T_5444 + _T_5445; // @[Bitwise.scala 48:55:@4862.4]
  assign _GEN_769 = {{1'd0}, _T_5443}; // @[Bitwise.scala 48:55:@4863.4]
  assign _T_5484 = _GEN_769 + _T_5483; // @[Bitwise.scala 48:55:@4863.4]
  assign _GEN_770 = {{1'd0}, _T_5482}; // @[Bitwise.scala 48:55:@4864.4]
  assign _T_5485 = _GEN_770 + _T_5484; // @[Bitwise.scala 48:55:@4864.4]
  assign _T_5486 = _T_5447 + _T_5448; // @[Bitwise.scala 48:55:@4865.4]
  assign _GEN_771 = {{1'd0}, _T_5446}; // @[Bitwise.scala 48:55:@4866.4]
  assign _T_5487 = _GEN_771 + _T_5486; // @[Bitwise.scala 48:55:@4866.4]
  assign _T_5488 = _T_5450 + _T_5451; // @[Bitwise.scala 48:55:@4867.4]
  assign _GEN_772 = {{1'd0}, _T_5449}; // @[Bitwise.scala 48:55:@4868.4]
  assign _T_5489 = _GEN_772 + _T_5488; // @[Bitwise.scala 48:55:@4868.4]
  assign _T_5490 = _T_5487 + _T_5489; // @[Bitwise.scala 48:55:@4869.4]
  assign _T_5491 = _T_5485 + _T_5490; // @[Bitwise.scala 48:55:@4870.4]
  assign _T_5492 = _T_5481 + _T_5491; // @[Bitwise.scala 48:55:@4871.4]
  assign _T_5493 = _T_5452 + _T_5453; // @[Bitwise.scala 48:55:@4872.4]
  assign _T_5494 = _T_5455 + _T_5456; // @[Bitwise.scala 48:55:@4873.4]
  assign _GEN_773 = {{1'd0}, _T_5454}; // @[Bitwise.scala 48:55:@4874.4]
  assign _T_5495 = _GEN_773 + _T_5494; // @[Bitwise.scala 48:55:@4874.4]
  assign _GEN_774 = {{1'd0}, _T_5493}; // @[Bitwise.scala 48:55:@4875.4]
  assign _T_5496 = _GEN_774 + _T_5495; // @[Bitwise.scala 48:55:@4875.4]
  assign _T_5497 = _T_5457 + _T_5458; // @[Bitwise.scala 48:55:@4876.4]
  assign _T_5498 = _T_5460 + _T_5461; // @[Bitwise.scala 48:55:@4877.4]
  assign _GEN_775 = {{1'd0}, _T_5459}; // @[Bitwise.scala 48:55:@4878.4]
  assign _T_5499 = _GEN_775 + _T_5498; // @[Bitwise.scala 48:55:@4878.4]
  assign _GEN_776 = {{1'd0}, _T_5497}; // @[Bitwise.scala 48:55:@4879.4]
  assign _T_5500 = _GEN_776 + _T_5499; // @[Bitwise.scala 48:55:@4879.4]
  assign _T_5501 = _T_5496 + _T_5500; // @[Bitwise.scala 48:55:@4880.4]
  assign _T_5502 = _T_5462 + _T_5463; // @[Bitwise.scala 48:55:@4881.4]
  assign _T_5503 = _T_5465 + _T_5466; // @[Bitwise.scala 48:55:@4882.4]
  assign _GEN_777 = {{1'd0}, _T_5464}; // @[Bitwise.scala 48:55:@4883.4]
  assign _T_5504 = _GEN_777 + _T_5503; // @[Bitwise.scala 48:55:@4883.4]
  assign _GEN_778 = {{1'd0}, _T_5502}; // @[Bitwise.scala 48:55:@4884.4]
  assign _T_5505 = _GEN_778 + _T_5504; // @[Bitwise.scala 48:55:@4884.4]
  assign _T_5506 = _T_5468 + _T_5469; // @[Bitwise.scala 48:55:@4885.4]
  assign _GEN_779 = {{1'd0}, _T_5467}; // @[Bitwise.scala 48:55:@4886.4]
  assign _T_5507 = _GEN_779 + _T_5506; // @[Bitwise.scala 48:55:@4886.4]
  assign _T_5508 = _T_5471 + _T_5472; // @[Bitwise.scala 48:55:@4887.4]
  assign _GEN_780 = {{1'd0}, _T_5470}; // @[Bitwise.scala 48:55:@4888.4]
  assign _T_5509 = _GEN_780 + _T_5508; // @[Bitwise.scala 48:55:@4888.4]
  assign _T_5510 = _T_5507 + _T_5509; // @[Bitwise.scala 48:55:@4889.4]
  assign _T_5511 = _T_5505 + _T_5510; // @[Bitwise.scala 48:55:@4890.4]
  assign _T_5512 = _T_5501 + _T_5511; // @[Bitwise.scala 48:55:@4891.4]
  assign _T_5513 = _T_5492 + _T_5512; // @[Bitwise.scala 48:55:@4892.4]
  assign _T_5577 = _T_1124[42:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@4957.4]
  assign _T_5578 = _T_5577[0]; // @[Bitwise.scala 50:65:@4958.4]
  assign _T_5579 = _T_5577[1]; // @[Bitwise.scala 50:65:@4959.4]
  assign _T_5580 = _T_5577[2]; // @[Bitwise.scala 50:65:@4960.4]
  assign _T_5581 = _T_5577[3]; // @[Bitwise.scala 50:65:@4961.4]
  assign _T_5582 = _T_5577[4]; // @[Bitwise.scala 50:65:@4962.4]
  assign _T_5583 = _T_5577[5]; // @[Bitwise.scala 50:65:@4963.4]
  assign _T_5584 = _T_5577[6]; // @[Bitwise.scala 50:65:@4964.4]
  assign _T_5585 = _T_5577[7]; // @[Bitwise.scala 50:65:@4965.4]
  assign _T_5586 = _T_5577[8]; // @[Bitwise.scala 50:65:@4966.4]
  assign _T_5587 = _T_5577[9]; // @[Bitwise.scala 50:65:@4967.4]
  assign _T_5588 = _T_5577[10]; // @[Bitwise.scala 50:65:@4968.4]
  assign _T_5589 = _T_5577[11]; // @[Bitwise.scala 50:65:@4969.4]
  assign _T_5590 = _T_5577[12]; // @[Bitwise.scala 50:65:@4970.4]
  assign _T_5591 = _T_5577[13]; // @[Bitwise.scala 50:65:@4971.4]
  assign _T_5592 = _T_5577[14]; // @[Bitwise.scala 50:65:@4972.4]
  assign _T_5593 = _T_5577[15]; // @[Bitwise.scala 50:65:@4973.4]
  assign _T_5594 = _T_5577[16]; // @[Bitwise.scala 50:65:@4974.4]
  assign _T_5595 = _T_5577[17]; // @[Bitwise.scala 50:65:@4975.4]
  assign _T_5596 = _T_5577[18]; // @[Bitwise.scala 50:65:@4976.4]
  assign _T_5597 = _T_5577[19]; // @[Bitwise.scala 50:65:@4977.4]
  assign _T_5598 = _T_5577[20]; // @[Bitwise.scala 50:65:@4978.4]
  assign _T_5599 = _T_5577[21]; // @[Bitwise.scala 50:65:@4979.4]
  assign _T_5600 = _T_5577[22]; // @[Bitwise.scala 50:65:@4980.4]
  assign _T_5601 = _T_5577[23]; // @[Bitwise.scala 50:65:@4981.4]
  assign _T_5602 = _T_5577[24]; // @[Bitwise.scala 50:65:@4982.4]
  assign _T_5603 = _T_5577[25]; // @[Bitwise.scala 50:65:@4983.4]
  assign _T_5604 = _T_5577[26]; // @[Bitwise.scala 50:65:@4984.4]
  assign _T_5605 = _T_5577[27]; // @[Bitwise.scala 50:65:@4985.4]
  assign _T_5606 = _T_5577[28]; // @[Bitwise.scala 50:65:@4986.4]
  assign _T_5607 = _T_5577[29]; // @[Bitwise.scala 50:65:@4987.4]
  assign _T_5608 = _T_5577[30]; // @[Bitwise.scala 50:65:@4988.4]
  assign _T_5609 = _T_5577[31]; // @[Bitwise.scala 50:65:@4989.4]
  assign _T_5610 = _T_5577[32]; // @[Bitwise.scala 50:65:@4990.4]
  assign _T_5611 = _T_5577[33]; // @[Bitwise.scala 50:65:@4991.4]
  assign _T_5612 = _T_5577[34]; // @[Bitwise.scala 50:65:@4992.4]
  assign _T_5613 = _T_5577[35]; // @[Bitwise.scala 50:65:@4993.4]
  assign _T_5614 = _T_5577[36]; // @[Bitwise.scala 50:65:@4994.4]
  assign _T_5615 = _T_5577[37]; // @[Bitwise.scala 50:65:@4995.4]
  assign _T_5616 = _T_5577[38]; // @[Bitwise.scala 50:65:@4996.4]
  assign _T_5617 = _T_5577[39]; // @[Bitwise.scala 50:65:@4997.4]
  assign _T_5618 = _T_5577[40]; // @[Bitwise.scala 50:65:@4998.4]
  assign _T_5619 = _T_5577[41]; // @[Bitwise.scala 50:65:@4999.4]
  assign _T_5620 = _T_5577[42]; // @[Bitwise.scala 50:65:@5000.4]
  assign _T_5621 = _T_5578 + _T_5579; // @[Bitwise.scala 48:55:@5001.4]
  assign _T_5622 = _T_5581 + _T_5582; // @[Bitwise.scala 48:55:@5002.4]
  assign _GEN_781 = {{1'd0}, _T_5580}; // @[Bitwise.scala 48:55:@5003.4]
  assign _T_5623 = _GEN_781 + _T_5622; // @[Bitwise.scala 48:55:@5003.4]
  assign _GEN_782 = {{1'd0}, _T_5621}; // @[Bitwise.scala 48:55:@5004.4]
  assign _T_5624 = _GEN_782 + _T_5623; // @[Bitwise.scala 48:55:@5004.4]
  assign _T_5625 = _T_5583 + _T_5584; // @[Bitwise.scala 48:55:@5005.4]
  assign _T_5626 = _T_5586 + _T_5587; // @[Bitwise.scala 48:55:@5006.4]
  assign _GEN_783 = {{1'd0}, _T_5585}; // @[Bitwise.scala 48:55:@5007.4]
  assign _T_5627 = _GEN_783 + _T_5626; // @[Bitwise.scala 48:55:@5007.4]
  assign _GEN_784 = {{1'd0}, _T_5625}; // @[Bitwise.scala 48:55:@5008.4]
  assign _T_5628 = _GEN_784 + _T_5627; // @[Bitwise.scala 48:55:@5008.4]
  assign _T_5629 = _T_5624 + _T_5628; // @[Bitwise.scala 48:55:@5009.4]
  assign _T_5630 = _T_5588 + _T_5589; // @[Bitwise.scala 48:55:@5010.4]
  assign _T_5631 = _T_5591 + _T_5592; // @[Bitwise.scala 48:55:@5011.4]
  assign _GEN_785 = {{1'd0}, _T_5590}; // @[Bitwise.scala 48:55:@5012.4]
  assign _T_5632 = _GEN_785 + _T_5631; // @[Bitwise.scala 48:55:@5012.4]
  assign _GEN_786 = {{1'd0}, _T_5630}; // @[Bitwise.scala 48:55:@5013.4]
  assign _T_5633 = _GEN_786 + _T_5632; // @[Bitwise.scala 48:55:@5013.4]
  assign _T_5634 = _T_5594 + _T_5595; // @[Bitwise.scala 48:55:@5014.4]
  assign _GEN_787 = {{1'd0}, _T_5593}; // @[Bitwise.scala 48:55:@5015.4]
  assign _T_5635 = _GEN_787 + _T_5634; // @[Bitwise.scala 48:55:@5015.4]
  assign _T_5636 = _T_5597 + _T_5598; // @[Bitwise.scala 48:55:@5016.4]
  assign _GEN_788 = {{1'd0}, _T_5596}; // @[Bitwise.scala 48:55:@5017.4]
  assign _T_5637 = _GEN_788 + _T_5636; // @[Bitwise.scala 48:55:@5017.4]
  assign _T_5638 = _T_5635 + _T_5637; // @[Bitwise.scala 48:55:@5018.4]
  assign _T_5639 = _T_5633 + _T_5638; // @[Bitwise.scala 48:55:@5019.4]
  assign _T_5640 = _T_5629 + _T_5639; // @[Bitwise.scala 48:55:@5020.4]
  assign _T_5641 = _T_5599 + _T_5600; // @[Bitwise.scala 48:55:@5021.4]
  assign _T_5642 = _T_5602 + _T_5603; // @[Bitwise.scala 48:55:@5022.4]
  assign _GEN_789 = {{1'd0}, _T_5601}; // @[Bitwise.scala 48:55:@5023.4]
  assign _T_5643 = _GEN_789 + _T_5642; // @[Bitwise.scala 48:55:@5023.4]
  assign _GEN_790 = {{1'd0}, _T_5641}; // @[Bitwise.scala 48:55:@5024.4]
  assign _T_5644 = _GEN_790 + _T_5643; // @[Bitwise.scala 48:55:@5024.4]
  assign _T_5645 = _T_5605 + _T_5606; // @[Bitwise.scala 48:55:@5025.4]
  assign _GEN_791 = {{1'd0}, _T_5604}; // @[Bitwise.scala 48:55:@5026.4]
  assign _T_5646 = _GEN_791 + _T_5645; // @[Bitwise.scala 48:55:@5026.4]
  assign _T_5647 = _T_5608 + _T_5609; // @[Bitwise.scala 48:55:@5027.4]
  assign _GEN_792 = {{1'd0}, _T_5607}; // @[Bitwise.scala 48:55:@5028.4]
  assign _T_5648 = _GEN_792 + _T_5647; // @[Bitwise.scala 48:55:@5028.4]
  assign _T_5649 = _T_5646 + _T_5648; // @[Bitwise.scala 48:55:@5029.4]
  assign _T_5650 = _T_5644 + _T_5649; // @[Bitwise.scala 48:55:@5030.4]
  assign _T_5651 = _T_5610 + _T_5611; // @[Bitwise.scala 48:55:@5031.4]
  assign _T_5652 = _T_5613 + _T_5614; // @[Bitwise.scala 48:55:@5032.4]
  assign _GEN_793 = {{1'd0}, _T_5612}; // @[Bitwise.scala 48:55:@5033.4]
  assign _T_5653 = _GEN_793 + _T_5652; // @[Bitwise.scala 48:55:@5033.4]
  assign _GEN_794 = {{1'd0}, _T_5651}; // @[Bitwise.scala 48:55:@5034.4]
  assign _T_5654 = _GEN_794 + _T_5653; // @[Bitwise.scala 48:55:@5034.4]
  assign _T_5655 = _T_5616 + _T_5617; // @[Bitwise.scala 48:55:@5035.4]
  assign _GEN_795 = {{1'd0}, _T_5615}; // @[Bitwise.scala 48:55:@5036.4]
  assign _T_5656 = _GEN_795 + _T_5655; // @[Bitwise.scala 48:55:@5036.4]
  assign _T_5657 = _T_5619 + _T_5620; // @[Bitwise.scala 48:55:@5037.4]
  assign _GEN_796 = {{1'd0}, _T_5618}; // @[Bitwise.scala 48:55:@5038.4]
  assign _T_5658 = _GEN_796 + _T_5657; // @[Bitwise.scala 48:55:@5038.4]
  assign _T_5659 = _T_5656 + _T_5658; // @[Bitwise.scala 48:55:@5039.4]
  assign _T_5660 = _T_5654 + _T_5659; // @[Bitwise.scala 48:55:@5040.4]
  assign _T_5661 = _T_5650 + _T_5660; // @[Bitwise.scala 48:55:@5041.4]
  assign _T_5662 = _T_5640 + _T_5661; // @[Bitwise.scala 48:55:@5042.4]
  assign _T_5726 = _T_1124[43:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5107.4]
  assign _T_5727 = _T_5726[0]; // @[Bitwise.scala 50:65:@5108.4]
  assign _T_5728 = _T_5726[1]; // @[Bitwise.scala 50:65:@5109.4]
  assign _T_5729 = _T_5726[2]; // @[Bitwise.scala 50:65:@5110.4]
  assign _T_5730 = _T_5726[3]; // @[Bitwise.scala 50:65:@5111.4]
  assign _T_5731 = _T_5726[4]; // @[Bitwise.scala 50:65:@5112.4]
  assign _T_5732 = _T_5726[5]; // @[Bitwise.scala 50:65:@5113.4]
  assign _T_5733 = _T_5726[6]; // @[Bitwise.scala 50:65:@5114.4]
  assign _T_5734 = _T_5726[7]; // @[Bitwise.scala 50:65:@5115.4]
  assign _T_5735 = _T_5726[8]; // @[Bitwise.scala 50:65:@5116.4]
  assign _T_5736 = _T_5726[9]; // @[Bitwise.scala 50:65:@5117.4]
  assign _T_5737 = _T_5726[10]; // @[Bitwise.scala 50:65:@5118.4]
  assign _T_5738 = _T_5726[11]; // @[Bitwise.scala 50:65:@5119.4]
  assign _T_5739 = _T_5726[12]; // @[Bitwise.scala 50:65:@5120.4]
  assign _T_5740 = _T_5726[13]; // @[Bitwise.scala 50:65:@5121.4]
  assign _T_5741 = _T_5726[14]; // @[Bitwise.scala 50:65:@5122.4]
  assign _T_5742 = _T_5726[15]; // @[Bitwise.scala 50:65:@5123.4]
  assign _T_5743 = _T_5726[16]; // @[Bitwise.scala 50:65:@5124.4]
  assign _T_5744 = _T_5726[17]; // @[Bitwise.scala 50:65:@5125.4]
  assign _T_5745 = _T_5726[18]; // @[Bitwise.scala 50:65:@5126.4]
  assign _T_5746 = _T_5726[19]; // @[Bitwise.scala 50:65:@5127.4]
  assign _T_5747 = _T_5726[20]; // @[Bitwise.scala 50:65:@5128.4]
  assign _T_5748 = _T_5726[21]; // @[Bitwise.scala 50:65:@5129.4]
  assign _T_5749 = _T_5726[22]; // @[Bitwise.scala 50:65:@5130.4]
  assign _T_5750 = _T_5726[23]; // @[Bitwise.scala 50:65:@5131.4]
  assign _T_5751 = _T_5726[24]; // @[Bitwise.scala 50:65:@5132.4]
  assign _T_5752 = _T_5726[25]; // @[Bitwise.scala 50:65:@5133.4]
  assign _T_5753 = _T_5726[26]; // @[Bitwise.scala 50:65:@5134.4]
  assign _T_5754 = _T_5726[27]; // @[Bitwise.scala 50:65:@5135.4]
  assign _T_5755 = _T_5726[28]; // @[Bitwise.scala 50:65:@5136.4]
  assign _T_5756 = _T_5726[29]; // @[Bitwise.scala 50:65:@5137.4]
  assign _T_5757 = _T_5726[30]; // @[Bitwise.scala 50:65:@5138.4]
  assign _T_5758 = _T_5726[31]; // @[Bitwise.scala 50:65:@5139.4]
  assign _T_5759 = _T_5726[32]; // @[Bitwise.scala 50:65:@5140.4]
  assign _T_5760 = _T_5726[33]; // @[Bitwise.scala 50:65:@5141.4]
  assign _T_5761 = _T_5726[34]; // @[Bitwise.scala 50:65:@5142.4]
  assign _T_5762 = _T_5726[35]; // @[Bitwise.scala 50:65:@5143.4]
  assign _T_5763 = _T_5726[36]; // @[Bitwise.scala 50:65:@5144.4]
  assign _T_5764 = _T_5726[37]; // @[Bitwise.scala 50:65:@5145.4]
  assign _T_5765 = _T_5726[38]; // @[Bitwise.scala 50:65:@5146.4]
  assign _T_5766 = _T_5726[39]; // @[Bitwise.scala 50:65:@5147.4]
  assign _T_5767 = _T_5726[40]; // @[Bitwise.scala 50:65:@5148.4]
  assign _T_5768 = _T_5726[41]; // @[Bitwise.scala 50:65:@5149.4]
  assign _T_5769 = _T_5726[42]; // @[Bitwise.scala 50:65:@5150.4]
  assign _T_5770 = _T_5726[43]; // @[Bitwise.scala 50:65:@5151.4]
  assign _T_5771 = _T_5727 + _T_5728; // @[Bitwise.scala 48:55:@5152.4]
  assign _T_5772 = _T_5730 + _T_5731; // @[Bitwise.scala 48:55:@5153.4]
  assign _GEN_797 = {{1'd0}, _T_5729}; // @[Bitwise.scala 48:55:@5154.4]
  assign _T_5773 = _GEN_797 + _T_5772; // @[Bitwise.scala 48:55:@5154.4]
  assign _GEN_798 = {{1'd0}, _T_5771}; // @[Bitwise.scala 48:55:@5155.4]
  assign _T_5774 = _GEN_798 + _T_5773; // @[Bitwise.scala 48:55:@5155.4]
  assign _T_5775 = _T_5733 + _T_5734; // @[Bitwise.scala 48:55:@5156.4]
  assign _GEN_799 = {{1'd0}, _T_5732}; // @[Bitwise.scala 48:55:@5157.4]
  assign _T_5776 = _GEN_799 + _T_5775; // @[Bitwise.scala 48:55:@5157.4]
  assign _T_5777 = _T_5736 + _T_5737; // @[Bitwise.scala 48:55:@5158.4]
  assign _GEN_800 = {{1'd0}, _T_5735}; // @[Bitwise.scala 48:55:@5159.4]
  assign _T_5778 = _GEN_800 + _T_5777; // @[Bitwise.scala 48:55:@5159.4]
  assign _T_5779 = _T_5776 + _T_5778; // @[Bitwise.scala 48:55:@5160.4]
  assign _T_5780 = _T_5774 + _T_5779; // @[Bitwise.scala 48:55:@5161.4]
  assign _T_5781 = _T_5738 + _T_5739; // @[Bitwise.scala 48:55:@5162.4]
  assign _T_5782 = _T_5741 + _T_5742; // @[Bitwise.scala 48:55:@5163.4]
  assign _GEN_801 = {{1'd0}, _T_5740}; // @[Bitwise.scala 48:55:@5164.4]
  assign _T_5783 = _GEN_801 + _T_5782; // @[Bitwise.scala 48:55:@5164.4]
  assign _GEN_802 = {{1'd0}, _T_5781}; // @[Bitwise.scala 48:55:@5165.4]
  assign _T_5784 = _GEN_802 + _T_5783; // @[Bitwise.scala 48:55:@5165.4]
  assign _T_5785 = _T_5744 + _T_5745; // @[Bitwise.scala 48:55:@5166.4]
  assign _GEN_803 = {{1'd0}, _T_5743}; // @[Bitwise.scala 48:55:@5167.4]
  assign _T_5786 = _GEN_803 + _T_5785; // @[Bitwise.scala 48:55:@5167.4]
  assign _T_5787 = _T_5747 + _T_5748; // @[Bitwise.scala 48:55:@5168.4]
  assign _GEN_804 = {{1'd0}, _T_5746}; // @[Bitwise.scala 48:55:@5169.4]
  assign _T_5788 = _GEN_804 + _T_5787; // @[Bitwise.scala 48:55:@5169.4]
  assign _T_5789 = _T_5786 + _T_5788; // @[Bitwise.scala 48:55:@5170.4]
  assign _T_5790 = _T_5784 + _T_5789; // @[Bitwise.scala 48:55:@5171.4]
  assign _T_5791 = _T_5780 + _T_5790; // @[Bitwise.scala 48:55:@5172.4]
  assign _T_5792 = _T_5749 + _T_5750; // @[Bitwise.scala 48:55:@5173.4]
  assign _T_5793 = _T_5752 + _T_5753; // @[Bitwise.scala 48:55:@5174.4]
  assign _GEN_805 = {{1'd0}, _T_5751}; // @[Bitwise.scala 48:55:@5175.4]
  assign _T_5794 = _GEN_805 + _T_5793; // @[Bitwise.scala 48:55:@5175.4]
  assign _GEN_806 = {{1'd0}, _T_5792}; // @[Bitwise.scala 48:55:@5176.4]
  assign _T_5795 = _GEN_806 + _T_5794; // @[Bitwise.scala 48:55:@5176.4]
  assign _T_5796 = _T_5755 + _T_5756; // @[Bitwise.scala 48:55:@5177.4]
  assign _GEN_807 = {{1'd0}, _T_5754}; // @[Bitwise.scala 48:55:@5178.4]
  assign _T_5797 = _GEN_807 + _T_5796; // @[Bitwise.scala 48:55:@5178.4]
  assign _T_5798 = _T_5758 + _T_5759; // @[Bitwise.scala 48:55:@5179.4]
  assign _GEN_808 = {{1'd0}, _T_5757}; // @[Bitwise.scala 48:55:@5180.4]
  assign _T_5799 = _GEN_808 + _T_5798; // @[Bitwise.scala 48:55:@5180.4]
  assign _T_5800 = _T_5797 + _T_5799; // @[Bitwise.scala 48:55:@5181.4]
  assign _T_5801 = _T_5795 + _T_5800; // @[Bitwise.scala 48:55:@5182.4]
  assign _T_5802 = _T_5760 + _T_5761; // @[Bitwise.scala 48:55:@5183.4]
  assign _T_5803 = _T_5763 + _T_5764; // @[Bitwise.scala 48:55:@5184.4]
  assign _GEN_809 = {{1'd0}, _T_5762}; // @[Bitwise.scala 48:55:@5185.4]
  assign _T_5804 = _GEN_809 + _T_5803; // @[Bitwise.scala 48:55:@5185.4]
  assign _GEN_810 = {{1'd0}, _T_5802}; // @[Bitwise.scala 48:55:@5186.4]
  assign _T_5805 = _GEN_810 + _T_5804; // @[Bitwise.scala 48:55:@5186.4]
  assign _T_5806 = _T_5766 + _T_5767; // @[Bitwise.scala 48:55:@5187.4]
  assign _GEN_811 = {{1'd0}, _T_5765}; // @[Bitwise.scala 48:55:@5188.4]
  assign _T_5807 = _GEN_811 + _T_5806; // @[Bitwise.scala 48:55:@5188.4]
  assign _T_5808 = _T_5769 + _T_5770; // @[Bitwise.scala 48:55:@5189.4]
  assign _GEN_812 = {{1'd0}, _T_5768}; // @[Bitwise.scala 48:55:@5190.4]
  assign _T_5809 = _GEN_812 + _T_5808; // @[Bitwise.scala 48:55:@5190.4]
  assign _T_5810 = _T_5807 + _T_5809; // @[Bitwise.scala 48:55:@5191.4]
  assign _T_5811 = _T_5805 + _T_5810; // @[Bitwise.scala 48:55:@5192.4]
  assign _T_5812 = _T_5801 + _T_5811; // @[Bitwise.scala 48:55:@5193.4]
  assign _T_5813 = _T_5791 + _T_5812; // @[Bitwise.scala 48:55:@5194.4]
  assign _T_5877 = _T_1124[44:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5259.4]
  assign _T_5878 = _T_5877[0]; // @[Bitwise.scala 50:65:@5260.4]
  assign _T_5879 = _T_5877[1]; // @[Bitwise.scala 50:65:@5261.4]
  assign _T_5880 = _T_5877[2]; // @[Bitwise.scala 50:65:@5262.4]
  assign _T_5881 = _T_5877[3]; // @[Bitwise.scala 50:65:@5263.4]
  assign _T_5882 = _T_5877[4]; // @[Bitwise.scala 50:65:@5264.4]
  assign _T_5883 = _T_5877[5]; // @[Bitwise.scala 50:65:@5265.4]
  assign _T_5884 = _T_5877[6]; // @[Bitwise.scala 50:65:@5266.4]
  assign _T_5885 = _T_5877[7]; // @[Bitwise.scala 50:65:@5267.4]
  assign _T_5886 = _T_5877[8]; // @[Bitwise.scala 50:65:@5268.4]
  assign _T_5887 = _T_5877[9]; // @[Bitwise.scala 50:65:@5269.4]
  assign _T_5888 = _T_5877[10]; // @[Bitwise.scala 50:65:@5270.4]
  assign _T_5889 = _T_5877[11]; // @[Bitwise.scala 50:65:@5271.4]
  assign _T_5890 = _T_5877[12]; // @[Bitwise.scala 50:65:@5272.4]
  assign _T_5891 = _T_5877[13]; // @[Bitwise.scala 50:65:@5273.4]
  assign _T_5892 = _T_5877[14]; // @[Bitwise.scala 50:65:@5274.4]
  assign _T_5893 = _T_5877[15]; // @[Bitwise.scala 50:65:@5275.4]
  assign _T_5894 = _T_5877[16]; // @[Bitwise.scala 50:65:@5276.4]
  assign _T_5895 = _T_5877[17]; // @[Bitwise.scala 50:65:@5277.4]
  assign _T_5896 = _T_5877[18]; // @[Bitwise.scala 50:65:@5278.4]
  assign _T_5897 = _T_5877[19]; // @[Bitwise.scala 50:65:@5279.4]
  assign _T_5898 = _T_5877[20]; // @[Bitwise.scala 50:65:@5280.4]
  assign _T_5899 = _T_5877[21]; // @[Bitwise.scala 50:65:@5281.4]
  assign _T_5900 = _T_5877[22]; // @[Bitwise.scala 50:65:@5282.4]
  assign _T_5901 = _T_5877[23]; // @[Bitwise.scala 50:65:@5283.4]
  assign _T_5902 = _T_5877[24]; // @[Bitwise.scala 50:65:@5284.4]
  assign _T_5903 = _T_5877[25]; // @[Bitwise.scala 50:65:@5285.4]
  assign _T_5904 = _T_5877[26]; // @[Bitwise.scala 50:65:@5286.4]
  assign _T_5905 = _T_5877[27]; // @[Bitwise.scala 50:65:@5287.4]
  assign _T_5906 = _T_5877[28]; // @[Bitwise.scala 50:65:@5288.4]
  assign _T_5907 = _T_5877[29]; // @[Bitwise.scala 50:65:@5289.4]
  assign _T_5908 = _T_5877[30]; // @[Bitwise.scala 50:65:@5290.4]
  assign _T_5909 = _T_5877[31]; // @[Bitwise.scala 50:65:@5291.4]
  assign _T_5910 = _T_5877[32]; // @[Bitwise.scala 50:65:@5292.4]
  assign _T_5911 = _T_5877[33]; // @[Bitwise.scala 50:65:@5293.4]
  assign _T_5912 = _T_5877[34]; // @[Bitwise.scala 50:65:@5294.4]
  assign _T_5913 = _T_5877[35]; // @[Bitwise.scala 50:65:@5295.4]
  assign _T_5914 = _T_5877[36]; // @[Bitwise.scala 50:65:@5296.4]
  assign _T_5915 = _T_5877[37]; // @[Bitwise.scala 50:65:@5297.4]
  assign _T_5916 = _T_5877[38]; // @[Bitwise.scala 50:65:@5298.4]
  assign _T_5917 = _T_5877[39]; // @[Bitwise.scala 50:65:@5299.4]
  assign _T_5918 = _T_5877[40]; // @[Bitwise.scala 50:65:@5300.4]
  assign _T_5919 = _T_5877[41]; // @[Bitwise.scala 50:65:@5301.4]
  assign _T_5920 = _T_5877[42]; // @[Bitwise.scala 50:65:@5302.4]
  assign _T_5921 = _T_5877[43]; // @[Bitwise.scala 50:65:@5303.4]
  assign _T_5922 = _T_5877[44]; // @[Bitwise.scala 50:65:@5304.4]
  assign _T_5923 = _T_5878 + _T_5879; // @[Bitwise.scala 48:55:@5305.4]
  assign _T_5924 = _T_5881 + _T_5882; // @[Bitwise.scala 48:55:@5306.4]
  assign _GEN_813 = {{1'd0}, _T_5880}; // @[Bitwise.scala 48:55:@5307.4]
  assign _T_5925 = _GEN_813 + _T_5924; // @[Bitwise.scala 48:55:@5307.4]
  assign _GEN_814 = {{1'd0}, _T_5923}; // @[Bitwise.scala 48:55:@5308.4]
  assign _T_5926 = _GEN_814 + _T_5925; // @[Bitwise.scala 48:55:@5308.4]
  assign _T_5927 = _T_5884 + _T_5885; // @[Bitwise.scala 48:55:@5309.4]
  assign _GEN_815 = {{1'd0}, _T_5883}; // @[Bitwise.scala 48:55:@5310.4]
  assign _T_5928 = _GEN_815 + _T_5927; // @[Bitwise.scala 48:55:@5310.4]
  assign _T_5929 = _T_5887 + _T_5888; // @[Bitwise.scala 48:55:@5311.4]
  assign _GEN_816 = {{1'd0}, _T_5886}; // @[Bitwise.scala 48:55:@5312.4]
  assign _T_5930 = _GEN_816 + _T_5929; // @[Bitwise.scala 48:55:@5312.4]
  assign _T_5931 = _T_5928 + _T_5930; // @[Bitwise.scala 48:55:@5313.4]
  assign _T_5932 = _T_5926 + _T_5931; // @[Bitwise.scala 48:55:@5314.4]
  assign _T_5933 = _T_5889 + _T_5890; // @[Bitwise.scala 48:55:@5315.4]
  assign _T_5934 = _T_5892 + _T_5893; // @[Bitwise.scala 48:55:@5316.4]
  assign _GEN_817 = {{1'd0}, _T_5891}; // @[Bitwise.scala 48:55:@5317.4]
  assign _T_5935 = _GEN_817 + _T_5934; // @[Bitwise.scala 48:55:@5317.4]
  assign _GEN_818 = {{1'd0}, _T_5933}; // @[Bitwise.scala 48:55:@5318.4]
  assign _T_5936 = _GEN_818 + _T_5935; // @[Bitwise.scala 48:55:@5318.4]
  assign _T_5937 = _T_5895 + _T_5896; // @[Bitwise.scala 48:55:@5319.4]
  assign _GEN_819 = {{1'd0}, _T_5894}; // @[Bitwise.scala 48:55:@5320.4]
  assign _T_5938 = _GEN_819 + _T_5937; // @[Bitwise.scala 48:55:@5320.4]
  assign _T_5939 = _T_5898 + _T_5899; // @[Bitwise.scala 48:55:@5321.4]
  assign _GEN_820 = {{1'd0}, _T_5897}; // @[Bitwise.scala 48:55:@5322.4]
  assign _T_5940 = _GEN_820 + _T_5939; // @[Bitwise.scala 48:55:@5322.4]
  assign _T_5941 = _T_5938 + _T_5940; // @[Bitwise.scala 48:55:@5323.4]
  assign _T_5942 = _T_5936 + _T_5941; // @[Bitwise.scala 48:55:@5324.4]
  assign _T_5943 = _T_5932 + _T_5942; // @[Bitwise.scala 48:55:@5325.4]
  assign _T_5944 = _T_5900 + _T_5901; // @[Bitwise.scala 48:55:@5326.4]
  assign _T_5945 = _T_5903 + _T_5904; // @[Bitwise.scala 48:55:@5327.4]
  assign _GEN_821 = {{1'd0}, _T_5902}; // @[Bitwise.scala 48:55:@5328.4]
  assign _T_5946 = _GEN_821 + _T_5945; // @[Bitwise.scala 48:55:@5328.4]
  assign _GEN_822 = {{1'd0}, _T_5944}; // @[Bitwise.scala 48:55:@5329.4]
  assign _T_5947 = _GEN_822 + _T_5946; // @[Bitwise.scala 48:55:@5329.4]
  assign _T_5948 = _T_5906 + _T_5907; // @[Bitwise.scala 48:55:@5330.4]
  assign _GEN_823 = {{1'd0}, _T_5905}; // @[Bitwise.scala 48:55:@5331.4]
  assign _T_5949 = _GEN_823 + _T_5948; // @[Bitwise.scala 48:55:@5331.4]
  assign _T_5950 = _T_5909 + _T_5910; // @[Bitwise.scala 48:55:@5332.4]
  assign _GEN_824 = {{1'd0}, _T_5908}; // @[Bitwise.scala 48:55:@5333.4]
  assign _T_5951 = _GEN_824 + _T_5950; // @[Bitwise.scala 48:55:@5333.4]
  assign _T_5952 = _T_5949 + _T_5951; // @[Bitwise.scala 48:55:@5334.4]
  assign _T_5953 = _T_5947 + _T_5952; // @[Bitwise.scala 48:55:@5335.4]
  assign _T_5954 = _T_5912 + _T_5913; // @[Bitwise.scala 48:55:@5336.4]
  assign _GEN_825 = {{1'd0}, _T_5911}; // @[Bitwise.scala 48:55:@5337.4]
  assign _T_5955 = _GEN_825 + _T_5954; // @[Bitwise.scala 48:55:@5337.4]
  assign _T_5956 = _T_5915 + _T_5916; // @[Bitwise.scala 48:55:@5338.4]
  assign _GEN_826 = {{1'd0}, _T_5914}; // @[Bitwise.scala 48:55:@5339.4]
  assign _T_5957 = _GEN_826 + _T_5956; // @[Bitwise.scala 48:55:@5339.4]
  assign _T_5958 = _T_5955 + _T_5957; // @[Bitwise.scala 48:55:@5340.4]
  assign _T_5959 = _T_5918 + _T_5919; // @[Bitwise.scala 48:55:@5341.4]
  assign _GEN_827 = {{1'd0}, _T_5917}; // @[Bitwise.scala 48:55:@5342.4]
  assign _T_5960 = _GEN_827 + _T_5959; // @[Bitwise.scala 48:55:@5342.4]
  assign _T_5961 = _T_5921 + _T_5922; // @[Bitwise.scala 48:55:@5343.4]
  assign _GEN_828 = {{1'd0}, _T_5920}; // @[Bitwise.scala 48:55:@5344.4]
  assign _T_5962 = _GEN_828 + _T_5961; // @[Bitwise.scala 48:55:@5344.4]
  assign _T_5963 = _T_5960 + _T_5962; // @[Bitwise.scala 48:55:@5345.4]
  assign _T_5964 = _T_5958 + _T_5963; // @[Bitwise.scala 48:55:@5346.4]
  assign _T_5965 = _T_5953 + _T_5964; // @[Bitwise.scala 48:55:@5347.4]
  assign _T_5966 = _T_5943 + _T_5965; // @[Bitwise.scala 48:55:@5348.4]
  assign _T_6030 = _T_1124[45:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5413.4]
  assign _T_6031 = _T_6030[0]; // @[Bitwise.scala 50:65:@5414.4]
  assign _T_6032 = _T_6030[1]; // @[Bitwise.scala 50:65:@5415.4]
  assign _T_6033 = _T_6030[2]; // @[Bitwise.scala 50:65:@5416.4]
  assign _T_6034 = _T_6030[3]; // @[Bitwise.scala 50:65:@5417.4]
  assign _T_6035 = _T_6030[4]; // @[Bitwise.scala 50:65:@5418.4]
  assign _T_6036 = _T_6030[5]; // @[Bitwise.scala 50:65:@5419.4]
  assign _T_6037 = _T_6030[6]; // @[Bitwise.scala 50:65:@5420.4]
  assign _T_6038 = _T_6030[7]; // @[Bitwise.scala 50:65:@5421.4]
  assign _T_6039 = _T_6030[8]; // @[Bitwise.scala 50:65:@5422.4]
  assign _T_6040 = _T_6030[9]; // @[Bitwise.scala 50:65:@5423.4]
  assign _T_6041 = _T_6030[10]; // @[Bitwise.scala 50:65:@5424.4]
  assign _T_6042 = _T_6030[11]; // @[Bitwise.scala 50:65:@5425.4]
  assign _T_6043 = _T_6030[12]; // @[Bitwise.scala 50:65:@5426.4]
  assign _T_6044 = _T_6030[13]; // @[Bitwise.scala 50:65:@5427.4]
  assign _T_6045 = _T_6030[14]; // @[Bitwise.scala 50:65:@5428.4]
  assign _T_6046 = _T_6030[15]; // @[Bitwise.scala 50:65:@5429.4]
  assign _T_6047 = _T_6030[16]; // @[Bitwise.scala 50:65:@5430.4]
  assign _T_6048 = _T_6030[17]; // @[Bitwise.scala 50:65:@5431.4]
  assign _T_6049 = _T_6030[18]; // @[Bitwise.scala 50:65:@5432.4]
  assign _T_6050 = _T_6030[19]; // @[Bitwise.scala 50:65:@5433.4]
  assign _T_6051 = _T_6030[20]; // @[Bitwise.scala 50:65:@5434.4]
  assign _T_6052 = _T_6030[21]; // @[Bitwise.scala 50:65:@5435.4]
  assign _T_6053 = _T_6030[22]; // @[Bitwise.scala 50:65:@5436.4]
  assign _T_6054 = _T_6030[23]; // @[Bitwise.scala 50:65:@5437.4]
  assign _T_6055 = _T_6030[24]; // @[Bitwise.scala 50:65:@5438.4]
  assign _T_6056 = _T_6030[25]; // @[Bitwise.scala 50:65:@5439.4]
  assign _T_6057 = _T_6030[26]; // @[Bitwise.scala 50:65:@5440.4]
  assign _T_6058 = _T_6030[27]; // @[Bitwise.scala 50:65:@5441.4]
  assign _T_6059 = _T_6030[28]; // @[Bitwise.scala 50:65:@5442.4]
  assign _T_6060 = _T_6030[29]; // @[Bitwise.scala 50:65:@5443.4]
  assign _T_6061 = _T_6030[30]; // @[Bitwise.scala 50:65:@5444.4]
  assign _T_6062 = _T_6030[31]; // @[Bitwise.scala 50:65:@5445.4]
  assign _T_6063 = _T_6030[32]; // @[Bitwise.scala 50:65:@5446.4]
  assign _T_6064 = _T_6030[33]; // @[Bitwise.scala 50:65:@5447.4]
  assign _T_6065 = _T_6030[34]; // @[Bitwise.scala 50:65:@5448.4]
  assign _T_6066 = _T_6030[35]; // @[Bitwise.scala 50:65:@5449.4]
  assign _T_6067 = _T_6030[36]; // @[Bitwise.scala 50:65:@5450.4]
  assign _T_6068 = _T_6030[37]; // @[Bitwise.scala 50:65:@5451.4]
  assign _T_6069 = _T_6030[38]; // @[Bitwise.scala 50:65:@5452.4]
  assign _T_6070 = _T_6030[39]; // @[Bitwise.scala 50:65:@5453.4]
  assign _T_6071 = _T_6030[40]; // @[Bitwise.scala 50:65:@5454.4]
  assign _T_6072 = _T_6030[41]; // @[Bitwise.scala 50:65:@5455.4]
  assign _T_6073 = _T_6030[42]; // @[Bitwise.scala 50:65:@5456.4]
  assign _T_6074 = _T_6030[43]; // @[Bitwise.scala 50:65:@5457.4]
  assign _T_6075 = _T_6030[44]; // @[Bitwise.scala 50:65:@5458.4]
  assign _T_6076 = _T_6030[45]; // @[Bitwise.scala 50:65:@5459.4]
  assign _T_6077 = _T_6031 + _T_6032; // @[Bitwise.scala 48:55:@5460.4]
  assign _T_6078 = _T_6034 + _T_6035; // @[Bitwise.scala 48:55:@5461.4]
  assign _GEN_829 = {{1'd0}, _T_6033}; // @[Bitwise.scala 48:55:@5462.4]
  assign _T_6079 = _GEN_829 + _T_6078; // @[Bitwise.scala 48:55:@5462.4]
  assign _GEN_830 = {{1'd0}, _T_6077}; // @[Bitwise.scala 48:55:@5463.4]
  assign _T_6080 = _GEN_830 + _T_6079; // @[Bitwise.scala 48:55:@5463.4]
  assign _T_6081 = _T_6037 + _T_6038; // @[Bitwise.scala 48:55:@5464.4]
  assign _GEN_831 = {{1'd0}, _T_6036}; // @[Bitwise.scala 48:55:@5465.4]
  assign _T_6082 = _GEN_831 + _T_6081; // @[Bitwise.scala 48:55:@5465.4]
  assign _T_6083 = _T_6040 + _T_6041; // @[Bitwise.scala 48:55:@5466.4]
  assign _GEN_832 = {{1'd0}, _T_6039}; // @[Bitwise.scala 48:55:@5467.4]
  assign _T_6084 = _GEN_832 + _T_6083; // @[Bitwise.scala 48:55:@5467.4]
  assign _T_6085 = _T_6082 + _T_6084; // @[Bitwise.scala 48:55:@5468.4]
  assign _T_6086 = _T_6080 + _T_6085; // @[Bitwise.scala 48:55:@5469.4]
  assign _T_6087 = _T_6043 + _T_6044; // @[Bitwise.scala 48:55:@5470.4]
  assign _GEN_833 = {{1'd0}, _T_6042}; // @[Bitwise.scala 48:55:@5471.4]
  assign _T_6088 = _GEN_833 + _T_6087; // @[Bitwise.scala 48:55:@5471.4]
  assign _T_6089 = _T_6046 + _T_6047; // @[Bitwise.scala 48:55:@5472.4]
  assign _GEN_834 = {{1'd0}, _T_6045}; // @[Bitwise.scala 48:55:@5473.4]
  assign _T_6090 = _GEN_834 + _T_6089; // @[Bitwise.scala 48:55:@5473.4]
  assign _T_6091 = _T_6088 + _T_6090; // @[Bitwise.scala 48:55:@5474.4]
  assign _T_6092 = _T_6049 + _T_6050; // @[Bitwise.scala 48:55:@5475.4]
  assign _GEN_835 = {{1'd0}, _T_6048}; // @[Bitwise.scala 48:55:@5476.4]
  assign _T_6093 = _GEN_835 + _T_6092; // @[Bitwise.scala 48:55:@5476.4]
  assign _T_6094 = _T_6052 + _T_6053; // @[Bitwise.scala 48:55:@5477.4]
  assign _GEN_836 = {{1'd0}, _T_6051}; // @[Bitwise.scala 48:55:@5478.4]
  assign _T_6095 = _GEN_836 + _T_6094; // @[Bitwise.scala 48:55:@5478.4]
  assign _T_6096 = _T_6093 + _T_6095; // @[Bitwise.scala 48:55:@5479.4]
  assign _T_6097 = _T_6091 + _T_6096; // @[Bitwise.scala 48:55:@5480.4]
  assign _T_6098 = _T_6086 + _T_6097; // @[Bitwise.scala 48:55:@5481.4]
  assign _T_6099 = _T_6054 + _T_6055; // @[Bitwise.scala 48:55:@5482.4]
  assign _T_6100 = _T_6057 + _T_6058; // @[Bitwise.scala 48:55:@5483.4]
  assign _GEN_837 = {{1'd0}, _T_6056}; // @[Bitwise.scala 48:55:@5484.4]
  assign _T_6101 = _GEN_837 + _T_6100; // @[Bitwise.scala 48:55:@5484.4]
  assign _GEN_838 = {{1'd0}, _T_6099}; // @[Bitwise.scala 48:55:@5485.4]
  assign _T_6102 = _GEN_838 + _T_6101; // @[Bitwise.scala 48:55:@5485.4]
  assign _T_6103 = _T_6060 + _T_6061; // @[Bitwise.scala 48:55:@5486.4]
  assign _GEN_839 = {{1'd0}, _T_6059}; // @[Bitwise.scala 48:55:@5487.4]
  assign _T_6104 = _GEN_839 + _T_6103; // @[Bitwise.scala 48:55:@5487.4]
  assign _T_6105 = _T_6063 + _T_6064; // @[Bitwise.scala 48:55:@5488.4]
  assign _GEN_840 = {{1'd0}, _T_6062}; // @[Bitwise.scala 48:55:@5489.4]
  assign _T_6106 = _GEN_840 + _T_6105; // @[Bitwise.scala 48:55:@5489.4]
  assign _T_6107 = _T_6104 + _T_6106; // @[Bitwise.scala 48:55:@5490.4]
  assign _T_6108 = _T_6102 + _T_6107; // @[Bitwise.scala 48:55:@5491.4]
  assign _T_6109 = _T_6066 + _T_6067; // @[Bitwise.scala 48:55:@5492.4]
  assign _GEN_841 = {{1'd0}, _T_6065}; // @[Bitwise.scala 48:55:@5493.4]
  assign _T_6110 = _GEN_841 + _T_6109; // @[Bitwise.scala 48:55:@5493.4]
  assign _T_6111 = _T_6069 + _T_6070; // @[Bitwise.scala 48:55:@5494.4]
  assign _GEN_842 = {{1'd0}, _T_6068}; // @[Bitwise.scala 48:55:@5495.4]
  assign _T_6112 = _GEN_842 + _T_6111; // @[Bitwise.scala 48:55:@5495.4]
  assign _T_6113 = _T_6110 + _T_6112; // @[Bitwise.scala 48:55:@5496.4]
  assign _T_6114 = _T_6072 + _T_6073; // @[Bitwise.scala 48:55:@5497.4]
  assign _GEN_843 = {{1'd0}, _T_6071}; // @[Bitwise.scala 48:55:@5498.4]
  assign _T_6115 = _GEN_843 + _T_6114; // @[Bitwise.scala 48:55:@5498.4]
  assign _T_6116 = _T_6075 + _T_6076; // @[Bitwise.scala 48:55:@5499.4]
  assign _GEN_844 = {{1'd0}, _T_6074}; // @[Bitwise.scala 48:55:@5500.4]
  assign _T_6117 = _GEN_844 + _T_6116; // @[Bitwise.scala 48:55:@5500.4]
  assign _T_6118 = _T_6115 + _T_6117; // @[Bitwise.scala 48:55:@5501.4]
  assign _T_6119 = _T_6113 + _T_6118; // @[Bitwise.scala 48:55:@5502.4]
  assign _T_6120 = _T_6108 + _T_6119; // @[Bitwise.scala 48:55:@5503.4]
  assign _T_6121 = _T_6098 + _T_6120; // @[Bitwise.scala 48:55:@5504.4]
  assign _T_6185 = _T_1124[46:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5569.4]
  assign _T_6186 = _T_6185[0]; // @[Bitwise.scala 50:65:@5570.4]
  assign _T_6187 = _T_6185[1]; // @[Bitwise.scala 50:65:@5571.4]
  assign _T_6188 = _T_6185[2]; // @[Bitwise.scala 50:65:@5572.4]
  assign _T_6189 = _T_6185[3]; // @[Bitwise.scala 50:65:@5573.4]
  assign _T_6190 = _T_6185[4]; // @[Bitwise.scala 50:65:@5574.4]
  assign _T_6191 = _T_6185[5]; // @[Bitwise.scala 50:65:@5575.4]
  assign _T_6192 = _T_6185[6]; // @[Bitwise.scala 50:65:@5576.4]
  assign _T_6193 = _T_6185[7]; // @[Bitwise.scala 50:65:@5577.4]
  assign _T_6194 = _T_6185[8]; // @[Bitwise.scala 50:65:@5578.4]
  assign _T_6195 = _T_6185[9]; // @[Bitwise.scala 50:65:@5579.4]
  assign _T_6196 = _T_6185[10]; // @[Bitwise.scala 50:65:@5580.4]
  assign _T_6197 = _T_6185[11]; // @[Bitwise.scala 50:65:@5581.4]
  assign _T_6198 = _T_6185[12]; // @[Bitwise.scala 50:65:@5582.4]
  assign _T_6199 = _T_6185[13]; // @[Bitwise.scala 50:65:@5583.4]
  assign _T_6200 = _T_6185[14]; // @[Bitwise.scala 50:65:@5584.4]
  assign _T_6201 = _T_6185[15]; // @[Bitwise.scala 50:65:@5585.4]
  assign _T_6202 = _T_6185[16]; // @[Bitwise.scala 50:65:@5586.4]
  assign _T_6203 = _T_6185[17]; // @[Bitwise.scala 50:65:@5587.4]
  assign _T_6204 = _T_6185[18]; // @[Bitwise.scala 50:65:@5588.4]
  assign _T_6205 = _T_6185[19]; // @[Bitwise.scala 50:65:@5589.4]
  assign _T_6206 = _T_6185[20]; // @[Bitwise.scala 50:65:@5590.4]
  assign _T_6207 = _T_6185[21]; // @[Bitwise.scala 50:65:@5591.4]
  assign _T_6208 = _T_6185[22]; // @[Bitwise.scala 50:65:@5592.4]
  assign _T_6209 = _T_6185[23]; // @[Bitwise.scala 50:65:@5593.4]
  assign _T_6210 = _T_6185[24]; // @[Bitwise.scala 50:65:@5594.4]
  assign _T_6211 = _T_6185[25]; // @[Bitwise.scala 50:65:@5595.4]
  assign _T_6212 = _T_6185[26]; // @[Bitwise.scala 50:65:@5596.4]
  assign _T_6213 = _T_6185[27]; // @[Bitwise.scala 50:65:@5597.4]
  assign _T_6214 = _T_6185[28]; // @[Bitwise.scala 50:65:@5598.4]
  assign _T_6215 = _T_6185[29]; // @[Bitwise.scala 50:65:@5599.4]
  assign _T_6216 = _T_6185[30]; // @[Bitwise.scala 50:65:@5600.4]
  assign _T_6217 = _T_6185[31]; // @[Bitwise.scala 50:65:@5601.4]
  assign _T_6218 = _T_6185[32]; // @[Bitwise.scala 50:65:@5602.4]
  assign _T_6219 = _T_6185[33]; // @[Bitwise.scala 50:65:@5603.4]
  assign _T_6220 = _T_6185[34]; // @[Bitwise.scala 50:65:@5604.4]
  assign _T_6221 = _T_6185[35]; // @[Bitwise.scala 50:65:@5605.4]
  assign _T_6222 = _T_6185[36]; // @[Bitwise.scala 50:65:@5606.4]
  assign _T_6223 = _T_6185[37]; // @[Bitwise.scala 50:65:@5607.4]
  assign _T_6224 = _T_6185[38]; // @[Bitwise.scala 50:65:@5608.4]
  assign _T_6225 = _T_6185[39]; // @[Bitwise.scala 50:65:@5609.4]
  assign _T_6226 = _T_6185[40]; // @[Bitwise.scala 50:65:@5610.4]
  assign _T_6227 = _T_6185[41]; // @[Bitwise.scala 50:65:@5611.4]
  assign _T_6228 = _T_6185[42]; // @[Bitwise.scala 50:65:@5612.4]
  assign _T_6229 = _T_6185[43]; // @[Bitwise.scala 50:65:@5613.4]
  assign _T_6230 = _T_6185[44]; // @[Bitwise.scala 50:65:@5614.4]
  assign _T_6231 = _T_6185[45]; // @[Bitwise.scala 50:65:@5615.4]
  assign _T_6232 = _T_6185[46]; // @[Bitwise.scala 50:65:@5616.4]
  assign _T_6233 = _T_6186 + _T_6187; // @[Bitwise.scala 48:55:@5617.4]
  assign _T_6234 = _T_6189 + _T_6190; // @[Bitwise.scala 48:55:@5618.4]
  assign _GEN_845 = {{1'd0}, _T_6188}; // @[Bitwise.scala 48:55:@5619.4]
  assign _T_6235 = _GEN_845 + _T_6234; // @[Bitwise.scala 48:55:@5619.4]
  assign _GEN_846 = {{1'd0}, _T_6233}; // @[Bitwise.scala 48:55:@5620.4]
  assign _T_6236 = _GEN_846 + _T_6235; // @[Bitwise.scala 48:55:@5620.4]
  assign _T_6237 = _T_6192 + _T_6193; // @[Bitwise.scala 48:55:@5621.4]
  assign _GEN_847 = {{1'd0}, _T_6191}; // @[Bitwise.scala 48:55:@5622.4]
  assign _T_6238 = _GEN_847 + _T_6237; // @[Bitwise.scala 48:55:@5622.4]
  assign _T_6239 = _T_6195 + _T_6196; // @[Bitwise.scala 48:55:@5623.4]
  assign _GEN_848 = {{1'd0}, _T_6194}; // @[Bitwise.scala 48:55:@5624.4]
  assign _T_6240 = _GEN_848 + _T_6239; // @[Bitwise.scala 48:55:@5624.4]
  assign _T_6241 = _T_6238 + _T_6240; // @[Bitwise.scala 48:55:@5625.4]
  assign _T_6242 = _T_6236 + _T_6241; // @[Bitwise.scala 48:55:@5626.4]
  assign _T_6243 = _T_6198 + _T_6199; // @[Bitwise.scala 48:55:@5627.4]
  assign _GEN_849 = {{1'd0}, _T_6197}; // @[Bitwise.scala 48:55:@5628.4]
  assign _T_6244 = _GEN_849 + _T_6243; // @[Bitwise.scala 48:55:@5628.4]
  assign _T_6245 = _T_6201 + _T_6202; // @[Bitwise.scala 48:55:@5629.4]
  assign _GEN_850 = {{1'd0}, _T_6200}; // @[Bitwise.scala 48:55:@5630.4]
  assign _T_6246 = _GEN_850 + _T_6245; // @[Bitwise.scala 48:55:@5630.4]
  assign _T_6247 = _T_6244 + _T_6246; // @[Bitwise.scala 48:55:@5631.4]
  assign _T_6248 = _T_6204 + _T_6205; // @[Bitwise.scala 48:55:@5632.4]
  assign _GEN_851 = {{1'd0}, _T_6203}; // @[Bitwise.scala 48:55:@5633.4]
  assign _T_6249 = _GEN_851 + _T_6248; // @[Bitwise.scala 48:55:@5633.4]
  assign _T_6250 = _T_6207 + _T_6208; // @[Bitwise.scala 48:55:@5634.4]
  assign _GEN_852 = {{1'd0}, _T_6206}; // @[Bitwise.scala 48:55:@5635.4]
  assign _T_6251 = _GEN_852 + _T_6250; // @[Bitwise.scala 48:55:@5635.4]
  assign _T_6252 = _T_6249 + _T_6251; // @[Bitwise.scala 48:55:@5636.4]
  assign _T_6253 = _T_6247 + _T_6252; // @[Bitwise.scala 48:55:@5637.4]
  assign _T_6254 = _T_6242 + _T_6253; // @[Bitwise.scala 48:55:@5638.4]
  assign _T_6255 = _T_6210 + _T_6211; // @[Bitwise.scala 48:55:@5639.4]
  assign _GEN_853 = {{1'd0}, _T_6209}; // @[Bitwise.scala 48:55:@5640.4]
  assign _T_6256 = _GEN_853 + _T_6255; // @[Bitwise.scala 48:55:@5640.4]
  assign _T_6257 = _T_6213 + _T_6214; // @[Bitwise.scala 48:55:@5641.4]
  assign _GEN_854 = {{1'd0}, _T_6212}; // @[Bitwise.scala 48:55:@5642.4]
  assign _T_6258 = _GEN_854 + _T_6257; // @[Bitwise.scala 48:55:@5642.4]
  assign _T_6259 = _T_6256 + _T_6258; // @[Bitwise.scala 48:55:@5643.4]
  assign _T_6260 = _T_6216 + _T_6217; // @[Bitwise.scala 48:55:@5644.4]
  assign _GEN_855 = {{1'd0}, _T_6215}; // @[Bitwise.scala 48:55:@5645.4]
  assign _T_6261 = _GEN_855 + _T_6260; // @[Bitwise.scala 48:55:@5645.4]
  assign _T_6262 = _T_6219 + _T_6220; // @[Bitwise.scala 48:55:@5646.4]
  assign _GEN_856 = {{1'd0}, _T_6218}; // @[Bitwise.scala 48:55:@5647.4]
  assign _T_6263 = _GEN_856 + _T_6262; // @[Bitwise.scala 48:55:@5647.4]
  assign _T_6264 = _T_6261 + _T_6263; // @[Bitwise.scala 48:55:@5648.4]
  assign _T_6265 = _T_6259 + _T_6264; // @[Bitwise.scala 48:55:@5649.4]
  assign _T_6266 = _T_6222 + _T_6223; // @[Bitwise.scala 48:55:@5650.4]
  assign _GEN_857 = {{1'd0}, _T_6221}; // @[Bitwise.scala 48:55:@5651.4]
  assign _T_6267 = _GEN_857 + _T_6266; // @[Bitwise.scala 48:55:@5651.4]
  assign _T_6268 = _T_6225 + _T_6226; // @[Bitwise.scala 48:55:@5652.4]
  assign _GEN_858 = {{1'd0}, _T_6224}; // @[Bitwise.scala 48:55:@5653.4]
  assign _T_6269 = _GEN_858 + _T_6268; // @[Bitwise.scala 48:55:@5653.4]
  assign _T_6270 = _T_6267 + _T_6269; // @[Bitwise.scala 48:55:@5654.4]
  assign _T_6271 = _T_6228 + _T_6229; // @[Bitwise.scala 48:55:@5655.4]
  assign _GEN_859 = {{1'd0}, _T_6227}; // @[Bitwise.scala 48:55:@5656.4]
  assign _T_6272 = _GEN_859 + _T_6271; // @[Bitwise.scala 48:55:@5656.4]
  assign _T_6273 = _T_6231 + _T_6232; // @[Bitwise.scala 48:55:@5657.4]
  assign _GEN_860 = {{1'd0}, _T_6230}; // @[Bitwise.scala 48:55:@5658.4]
  assign _T_6274 = _GEN_860 + _T_6273; // @[Bitwise.scala 48:55:@5658.4]
  assign _T_6275 = _T_6272 + _T_6274; // @[Bitwise.scala 48:55:@5659.4]
  assign _T_6276 = _T_6270 + _T_6275; // @[Bitwise.scala 48:55:@5660.4]
  assign _T_6277 = _T_6265 + _T_6276; // @[Bitwise.scala 48:55:@5661.4]
  assign _T_6278 = _T_6254 + _T_6277; // @[Bitwise.scala 48:55:@5662.4]
  assign _T_6342 = _T_1124[47:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5727.4]
  assign _T_6343 = _T_6342[0]; // @[Bitwise.scala 50:65:@5728.4]
  assign _T_6344 = _T_6342[1]; // @[Bitwise.scala 50:65:@5729.4]
  assign _T_6345 = _T_6342[2]; // @[Bitwise.scala 50:65:@5730.4]
  assign _T_6346 = _T_6342[3]; // @[Bitwise.scala 50:65:@5731.4]
  assign _T_6347 = _T_6342[4]; // @[Bitwise.scala 50:65:@5732.4]
  assign _T_6348 = _T_6342[5]; // @[Bitwise.scala 50:65:@5733.4]
  assign _T_6349 = _T_6342[6]; // @[Bitwise.scala 50:65:@5734.4]
  assign _T_6350 = _T_6342[7]; // @[Bitwise.scala 50:65:@5735.4]
  assign _T_6351 = _T_6342[8]; // @[Bitwise.scala 50:65:@5736.4]
  assign _T_6352 = _T_6342[9]; // @[Bitwise.scala 50:65:@5737.4]
  assign _T_6353 = _T_6342[10]; // @[Bitwise.scala 50:65:@5738.4]
  assign _T_6354 = _T_6342[11]; // @[Bitwise.scala 50:65:@5739.4]
  assign _T_6355 = _T_6342[12]; // @[Bitwise.scala 50:65:@5740.4]
  assign _T_6356 = _T_6342[13]; // @[Bitwise.scala 50:65:@5741.4]
  assign _T_6357 = _T_6342[14]; // @[Bitwise.scala 50:65:@5742.4]
  assign _T_6358 = _T_6342[15]; // @[Bitwise.scala 50:65:@5743.4]
  assign _T_6359 = _T_6342[16]; // @[Bitwise.scala 50:65:@5744.4]
  assign _T_6360 = _T_6342[17]; // @[Bitwise.scala 50:65:@5745.4]
  assign _T_6361 = _T_6342[18]; // @[Bitwise.scala 50:65:@5746.4]
  assign _T_6362 = _T_6342[19]; // @[Bitwise.scala 50:65:@5747.4]
  assign _T_6363 = _T_6342[20]; // @[Bitwise.scala 50:65:@5748.4]
  assign _T_6364 = _T_6342[21]; // @[Bitwise.scala 50:65:@5749.4]
  assign _T_6365 = _T_6342[22]; // @[Bitwise.scala 50:65:@5750.4]
  assign _T_6366 = _T_6342[23]; // @[Bitwise.scala 50:65:@5751.4]
  assign _T_6367 = _T_6342[24]; // @[Bitwise.scala 50:65:@5752.4]
  assign _T_6368 = _T_6342[25]; // @[Bitwise.scala 50:65:@5753.4]
  assign _T_6369 = _T_6342[26]; // @[Bitwise.scala 50:65:@5754.4]
  assign _T_6370 = _T_6342[27]; // @[Bitwise.scala 50:65:@5755.4]
  assign _T_6371 = _T_6342[28]; // @[Bitwise.scala 50:65:@5756.4]
  assign _T_6372 = _T_6342[29]; // @[Bitwise.scala 50:65:@5757.4]
  assign _T_6373 = _T_6342[30]; // @[Bitwise.scala 50:65:@5758.4]
  assign _T_6374 = _T_6342[31]; // @[Bitwise.scala 50:65:@5759.4]
  assign _T_6375 = _T_6342[32]; // @[Bitwise.scala 50:65:@5760.4]
  assign _T_6376 = _T_6342[33]; // @[Bitwise.scala 50:65:@5761.4]
  assign _T_6377 = _T_6342[34]; // @[Bitwise.scala 50:65:@5762.4]
  assign _T_6378 = _T_6342[35]; // @[Bitwise.scala 50:65:@5763.4]
  assign _T_6379 = _T_6342[36]; // @[Bitwise.scala 50:65:@5764.4]
  assign _T_6380 = _T_6342[37]; // @[Bitwise.scala 50:65:@5765.4]
  assign _T_6381 = _T_6342[38]; // @[Bitwise.scala 50:65:@5766.4]
  assign _T_6382 = _T_6342[39]; // @[Bitwise.scala 50:65:@5767.4]
  assign _T_6383 = _T_6342[40]; // @[Bitwise.scala 50:65:@5768.4]
  assign _T_6384 = _T_6342[41]; // @[Bitwise.scala 50:65:@5769.4]
  assign _T_6385 = _T_6342[42]; // @[Bitwise.scala 50:65:@5770.4]
  assign _T_6386 = _T_6342[43]; // @[Bitwise.scala 50:65:@5771.4]
  assign _T_6387 = _T_6342[44]; // @[Bitwise.scala 50:65:@5772.4]
  assign _T_6388 = _T_6342[45]; // @[Bitwise.scala 50:65:@5773.4]
  assign _T_6389 = _T_6342[46]; // @[Bitwise.scala 50:65:@5774.4]
  assign _T_6390 = _T_6342[47]; // @[Bitwise.scala 50:65:@5775.4]
  assign _T_6391 = _T_6344 + _T_6345; // @[Bitwise.scala 48:55:@5776.4]
  assign _GEN_861 = {{1'd0}, _T_6343}; // @[Bitwise.scala 48:55:@5777.4]
  assign _T_6392 = _GEN_861 + _T_6391; // @[Bitwise.scala 48:55:@5777.4]
  assign _T_6393 = _T_6347 + _T_6348; // @[Bitwise.scala 48:55:@5778.4]
  assign _GEN_862 = {{1'd0}, _T_6346}; // @[Bitwise.scala 48:55:@5779.4]
  assign _T_6394 = _GEN_862 + _T_6393; // @[Bitwise.scala 48:55:@5779.4]
  assign _T_6395 = _T_6392 + _T_6394; // @[Bitwise.scala 48:55:@5780.4]
  assign _T_6396 = _T_6350 + _T_6351; // @[Bitwise.scala 48:55:@5781.4]
  assign _GEN_863 = {{1'd0}, _T_6349}; // @[Bitwise.scala 48:55:@5782.4]
  assign _T_6397 = _GEN_863 + _T_6396; // @[Bitwise.scala 48:55:@5782.4]
  assign _T_6398 = _T_6353 + _T_6354; // @[Bitwise.scala 48:55:@5783.4]
  assign _GEN_864 = {{1'd0}, _T_6352}; // @[Bitwise.scala 48:55:@5784.4]
  assign _T_6399 = _GEN_864 + _T_6398; // @[Bitwise.scala 48:55:@5784.4]
  assign _T_6400 = _T_6397 + _T_6399; // @[Bitwise.scala 48:55:@5785.4]
  assign _T_6401 = _T_6395 + _T_6400; // @[Bitwise.scala 48:55:@5786.4]
  assign _T_6402 = _T_6356 + _T_6357; // @[Bitwise.scala 48:55:@5787.4]
  assign _GEN_865 = {{1'd0}, _T_6355}; // @[Bitwise.scala 48:55:@5788.4]
  assign _T_6403 = _GEN_865 + _T_6402; // @[Bitwise.scala 48:55:@5788.4]
  assign _T_6404 = _T_6359 + _T_6360; // @[Bitwise.scala 48:55:@5789.4]
  assign _GEN_866 = {{1'd0}, _T_6358}; // @[Bitwise.scala 48:55:@5790.4]
  assign _T_6405 = _GEN_866 + _T_6404; // @[Bitwise.scala 48:55:@5790.4]
  assign _T_6406 = _T_6403 + _T_6405; // @[Bitwise.scala 48:55:@5791.4]
  assign _T_6407 = _T_6362 + _T_6363; // @[Bitwise.scala 48:55:@5792.4]
  assign _GEN_867 = {{1'd0}, _T_6361}; // @[Bitwise.scala 48:55:@5793.4]
  assign _T_6408 = _GEN_867 + _T_6407; // @[Bitwise.scala 48:55:@5793.4]
  assign _T_6409 = _T_6365 + _T_6366; // @[Bitwise.scala 48:55:@5794.4]
  assign _GEN_868 = {{1'd0}, _T_6364}; // @[Bitwise.scala 48:55:@5795.4]
  assign _T_6410 = _GEN_868 + _T_6409; // @[Bitwise.scala 48:55:@5795.4]
  assign _T_6411 = _T_6408 + _T_6410; // @[Bitwise.scala 48:55:@5796.4]
  assign _T_6412 = _T_6406 + _T_6411; // @[Bitwise.scala 48:55:@5797.4]
  assign _T_6413 = _T_6401 + _T_6412; // @[Bitwise.scala 48:55:@5798.4]
  assign _T_6414 = _T_6368 + _T_6369; // @[Bitwise.scala 48:55:@5799.4]
  assign _GEN_869 = {{1'd0}, _T_6367}; // @[Bitwise.scala 48:55:@5800.4]
  assign _T_6415 = _GEN_869 + _T_6414; // @[Bitwise.scala 48:55:@5800.4]
  assign _T_6416 = _T_6371 + _T_6372; // @[Bitwise.scala 48:55:@5801.4]
  assign _GEN_870 = {{1'd0}, _T_6370}; // @[Bitwise.scala 48:55:@5802.4]
  assign _T_6417 = _GEN_870 + _T_6416; // @[Bitwise.scala 48:55:@5802.4]
  assign _T_6418 = _T_6415 + _T_6417; // @[Bitwise.scala 48:55:@5803.4]
  assign _T_6419 = _T_6374 + _T_6375; // @[Bitwise.scala 48:55:@5804.4]
  assign _GEN_871 = {{1'd0}, _T_6373}; // @[Bitwise.scala 48:55:@5805.4]
  assign _T_6420 = _GEN_871 + _T_6419; // @[Bitwise.scala 48:55:@5805.4]
  assign _T_6421 = _T_6377 + _T_6378; // @[Bitwise.scala 48:55:@5806.4]
  assign _GEN_872 = {{1'd0}, _T_6376}; // @[Bitwise.scala 48:55:@5807.4]
  assign _T_6422 = _GEN_872 + _T_6421; // @[Bitwise.scala 48:55:@5807.4]
  assign _T_6423 = _T_6420 + _T_6422; // @[Bitwise.scala 48:55:@5808.4]
  assign _T_6424 = _T_6418 + _T_6423; // @[Bitwise.scala 48:55:@5809.4]
  assign _T_6425 = _T_6380 + _T_6381; // @[Bitwise.scala 48:55:@5810.4]
  assign _GEN_873 = {{1'd0}, _T_6379}; // @[Bitwise.scala 48:55:@5811.4]
  assign _T_6426 = _GEN_873 + _T_6425; // @[Bitwise.scala 48:55:@5811.4]
  assign _T_6427 = _T_6383 + _T_6384; // @[Bitwise.scala 48:55:@5812.4]
  assign _GEN_874 = {{1'd0}, _T_6382}; // @[Bitwise.scala 48:55:@5813.4]
  assign _T_6428 = _GEN_874 + _T_6427; // @[Bitwise.scala 48:55:@5813.4]
  assign _T_6429 = _T_6426 + _T_6428; // @[Bitwise.scala 48:55:@5814.4]
  assign _T_6430 = _T_6386 + _T_6387; // @[Bitwise.scala 48:55:@5815.4]
  assign _GEN_875 = {{1'd0}, _T_6385}; // @[Bitwise.scala 48:55:@5816.4]
  assign _T_6431 = _GEN_875 + _T_6430; // @[Bitwise.scala 48:55:@5816.4]
  assign _T_6432 = _T_6389 + _T_6390; // @[Bitwise.scala 48:55:@5817.4]
  assign _GEN_876 = {{1'd0}, _T_6388}; // @[Bitwise.scala 48:55:@5818.4]
  assign _T_6433 = _GEN_876 + _T_6432; // @[Bitwise.scala 48:55:@5818.4]
  assign _T_6434 = _T_6431 + _T_6433; // @[Bitwise.scala 48:55:@5819.4]
  assign _T_6435 = _T_6429 + _T_6434; // @[Bitwise.scala 48:55:@5820.4]
  assign _T_6436 = _T_6424 + _T_6435; // @[Bitwise.scala 48:55:@5821.4]
  assign _T_6437 = _T_6413 + _T_6436; // @[Bitwise.scala 48:55:@5822.4]
  assign _T_6501 = _T_1124[48:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@5887.4]
  assign _T_6502 = _T_6501[0]; // @[Bitwise.scala 50:65:@5888.4]
  assign _T_6503 = _T_6501[1]; // @[Bitwise.scala 50:65:@5889.4]
  assign _T_6504 = _T_6501[2]; // @[Bitwise.scala 50:65:@5890.4]
  assign _T_6505 = _T_6501[3]; // @[Bitwise.scala 50:65:@5891.4]
  assign _T_6506 = _T_6501[4]; // @[Bitwise.scala 50:65:@5892.4]
  assign _T_6507 = _T_6501[5]; // @[Bitwise.scala 50:65:@5893.4]
  assign _T_6508 = _T_6501[6]; // @[Bitwise.scala 50:65:@5894.4]
  assign _T_6509 = _T_6501[7]; // @[Bitwise.scala 50:65:@5895.4]
  assign _T_6510 = _T_6501[8]; // @[Bitwise.scala 50:65:@5896.4]
  assign _T_6511 = _T_6501[9]; // @[Bitwise.scala 50:65:@5897.4]
  assign _T_6512 = _T_6501[10]; // @[Bitwise.scala 50:65:@5898.4]
  assign _T_6513 = _T_6501[11]; // @[Bitwise.scala 50:65:@5899.4]
  assign _T_6514 = _T_6501[12]; // @[Bitwise.scala 50:65:@5900.4]
  assign _T_6515 = _T_6501[13]; // @[Bitwise.scala 50:65:@5901.4]
  assign _T_6516 = _T_6501[14]; // @[Bitwise.scala 50:65:@5902.4]
  assign _T_6517 = _T_6501[15]; // @[Bitwise.scala 50:65:@5903.4]
  assign _T_6518 = _T_6501[16]; // @[Bitwise.scala 50:65:@5904.4]
  assign _T_6519 = _T_6501[17]; // @[Bitwise.scala 50:65:@5905.4]
  assign _T_6520 = _T_6501[18]; // @[Bitwise.scala 50:65:@5906.4]
  assign _T_6521 = _T_6501[19]; // @[Bitwise.scala 50:65:@5907.4]
  assign _T_6522 = _T_6501[20]; // @[Bitwise.scala 50:65:@5908.4]
  assign _T_6523 = _T_6501[21]; // @[Bitwise.scala 50:65:@5909.4]
  assign _T_6524 = _T_6501[22]; // @[Bitwise.scala 50:65:@5910.4]
  assign _T_6525 = _T_6501[23]; // @[Bitwise.scala 50:65:@5911.4]
  assign _T_6526 = _T_6501[24]; // @[Bitwise.scala 50:65:@5912.4]
  assign _T_6527 = _T_6501[25]; // @[Bitwise.scala 50:65:@5913.4]
  assign _T_6528 = _T_6501[26]; // @[Bitwise.scala 50:65:@5914.4]
  assign _T_6529 = _T_6501[27]; // @[Bitwise.scala 50:65:@5915.4]
  assign _T_6530 = _T_6501[28]; // @[Bitwise.scala 50:65:@5916.4]
  assign _T_6531 = _T_6501[29]; // @[Bitwise.scala 50:65:@5917.4]
  assign _T_6532 = _T_6501[30]; // @[Bitwise.scala 50:65:@5918.4]
  assign _T_6533 = _T_6501[31]; // @[Bitwise.scala 50:65:@5919.4]
  assign _T_6534 = _T_6501[32]; // @[Bitwise.scala 50:65:@5920.4]
  assign _T_6535 = _T_6501[33]; // @[Bitwise.scala 50:65:@5921.4]
  assign _T_6536 = _T_6501[34]; // @[Bitwise.scala 50:65:@5922.4]
  assign _T_6537 = _T_6501[35]; // @[Bitwise.scala 50:65:@5923.4]
  assign _T_6538 = _T_6501[36]; // @[Bitwise.scala 50:65:@5924.4]
  assign _T_6539 = _T_6501[37]; // @[Bitwise.scala 50:65:@5925.4]
  assign _T_6540 = _T_6501[38]; // @[Bitwise.scala 50:65:@5926.4]
  assign _T_6541 = _T_6501[39]; // @[Bitwise.scala 50:65:@5927.4]
  assign _T_6542 = _T_6501[40]; // @[Bitwise.scala 50:65:@5928.4]
  assign _T_6543 = _T_6501[41]; // @[Bitwise.scala 50:65:@5929.4]
  assign _T_6544 = _T_6501[42]; // @[Bitwise.scala 50:65:@5930.4]
  assign _T_6545 = _T_6501[43]; // @[Bitwise.scala 50:65:@5931.4]
  assign _T_6546 = _T_6501[44]; // @[Bitwise.scala 50:65:@5932.4]
  assign _T_6547 = _T_6501[45]; // @[Bitwise.scala 50:65:@5933.4]
  assign _T_6548 = _T_6501[46]; // @[Bitwise.scala 50:65:@5934.4]
  assign _T_6549 = _T_6501[47]; // @[Bitwise.scala 50:65:@5935.4]
  assign _T_6550 = _T_6501[48]; // @[Bitwise.scala 50:65:@5936.4]
  assign _T_6551 = _T_6503 + _T_6504; // @[Bitwise.scala 48:55:@5937.4]
  assign _GEN_877 = {{1'd0}, _T_6502}; // @[Bitwise.scala 48:55:@5938.4]
  assign _T_6552 = _GEN_877 + _T_6551; // @[Bitwise.scala 48:55:@5938.4]
  assign _T_6553 = _T_6506 + _T_6507; // @[Bitwise.scala 48:55:@5939.4]
  assign _GEN_878 = {{1'd0}, _T_6505}; // @[Bitwise.scala 48:55:@5940.4]
  assign _T_6554 = _GEN_878 + _T_6553; // @[Bitwise.scala 48:55:@5940.4]
  assign _T_6555 = _T_6552 + _T_6554; // @[Bitwise.scala 48:55:@5941.4]
  assign _T_6556 = _T_6509 + _T_6510; // @[Bitwise.scala 48:55:@5942.4]
  assign _GEN_879 = {{1'd0}, _T_6508}; // @[Bitwise.scala 48:55:@5943.4]
  assign _T_6557 = _GEN_879 + _T_6556; // @[Bitwise.scala 48:55:@5943.4]
  assign _T_6558 = _T_6512 + _T_6513; // @[Bitwise.scala 48:55:@5944.4]
  assign _GEN_880 = {{1'd0}, _T_6511}; // @[Bitwise.scala 48:55:@5945.4]
  assign _T_6559 = _GEN_880 + _T_6558; // @[Bitwise.scala 48:55:@5945.4]
  assign _T_6560 = _T_6557 + _T_6559; // @[Bitwise.scala 48:55:@5946.4]
  assign _T_6561 = _T_6555 + _T_6560; // @[Bitwise.scala 48:55:@5947.4]
  assign _T_6562 = _T_6515 + _T_6516; // @[Bitwise.scala 48:55:@5948.4]
  assign _GEN_881 = {{1'd0}, _T_6514}; // @[Bitwise.scala 48:55:@5949.4]
  assign _T_6563 = _GEN_881 + _T_6562; // @[Bitwise.scala 48:55:@5949.4]
  assign _T_6564 = _T_6518 + _T_6519; // @[Bitwise.scala 48:55:@5950.4]
  assign _GEN_882 = {{1'd0}, _T_6517}; // @[Bitwise.scala 48:55:@5951.4]
  assign _T_6565 = _GEN_882 + _T_6564; // @[Bitwise.scala 48:55:@5951.4]
  assign _T_6566 = _T_6563 + _T_6565; // @[Bitwise.scala 48:55:@5952.4]
  assign _T_6567 = _T_6521 + _T_6522; // @[Bitwise.scala 48:55:@5953.4]
  assign _GEN_883 = {{1'd0}, _T_6520}; // @[Bitwise.scala 48:55:@5954.4]
  assign _T_6568 = _GEN_883 + _T_6567; // @[Bitwise.scala 48:55:@5954.4]
  assign _T_6569 = _T_6524 + _T_6525; // @[Bitwise.scala 48:55:@5955.4]
  assign _GEN_884 = {{1'd0}, _T_6523}; // @[Bitwise.scala 48:55:@5956.4]
  assign _T_6570 = _GEN_884 + _T_6569; // @[Bitwise.scala 48:55:@5956.4]
  assign _T_6571 = _T_6568 + _T_6570; // @[Bitwise.scala 48:55:@5957.4]
  assign _T_6572 = _T_6566 + _T_6571; // @[Bitwise.scala 48:55:@5958.4]
  assign _T_6573 = _T_6561 + _T_6572; // @[Bitwise.scala 48:55:@5959.4]
  assign _T_6574 = _T_6527 + _T_6528; // @[Bitwise.scala 48:55:@5960.4]
  assign _GEN_885 = {{1'd0}, _T_6526}; // @[Bitwise.scala 48:55:@5961.4]
  assign _T_6575 = _GEN_885 + _T_6574; // @[Bitwise.scala 48:55:@5961.4]
  assign _T_6576 = _T_6530 + _T_6531; // @[Bitwise.scala 48:55:@5962.4]
  assign _GEN_886 = {{1'd0}, _T_6529}; // @[Bitwise.scala 48:55:@5963.4]
  assign _T_6577 = _GEN_886 + _T_6576; // @[Bitwise.scala 48:55:@5963.4]
  assign _T_6578 = _T_6575 + _T_6577; // @[Bitwise.scala 48:55:@5964.4]
  assign _T_6579 = _T_6533 + _T_6534; // @[Bitwise.scala 48:55:@5965.4]
  assign _GEN_887 = {{1'd0}, _T_6532}; // @[Bitwise.scala 48:55:@5966.4]
  assign _T_6580 = _GEN_887 + _T_6579; // @[Bitwise.scala 48:55:@5966.4]
  assign _T_6581 = _T_6536 + _T_6537; // @[Bitwise.scala 48:55:@5967.4]
  assign _GEN_888 = {{1'd0}, _T_6535}; // @[Bitwise.scala 48:55:@5968.4]
  assign _T_6582 = _GEN_888 + _T_6581; // @[Bitwise.scala 48:55:@5968.4]
  assign _T_6583 = _T_6580 + _T_6582; // @[Bitwise.scala 48:55:@5969.4]
  assign _T_6584 = _T_6578 + _T_6583; // @[Bitwise.scala 48:55:@5970.4]
  assign _T_6585 = _T_6539 + _T_6540; // @[Bitwise.scala 48:55:@5971.4]
  assign _GEN_889 = {{1'd0}, _T_6538}; // @[Bitwise.scala 48:55:@5972.4]
  assign _T_6586 = _GEN_889 + _T_6585; // @[Bitwise.scala 48:55:@5972.4]
  assign _T_6587 = _T_6542 + _T_6543; // @[Bitwise.scala 48:55:@5973.4]
  assign _GEN_890 = {{1'd0}, _T_6541}; // @[Bitwise.scala 48:55:@5974.4]
  assign _T_6588 = _GEN_890 + _T_6587; // @[Bitwise.scala 48:55:@5974.4]
  assign _T_6589 = _T_6586 + _T_6588; // @[Bitwise.scala 48:55:@5975.4]
  assign _T_6590 = _T_6545 + _T_6546; // @[Bitwise.scala 48:55:@5976.4]
  assign _GEN_891 = {{1'd0}, _T_6544}; // @[Bitwise.scala 48:55:@5977.4]
  assign _T_6591 = _GEN_891 + _T_6590; // @[Bitwise.scala 48:55:@5977.4]
  assign _T_6592 = _T_6547 + _T_6548; // @[Bitwise.scala 48:55:@5978.4]
  assign _T_6593 = _T_6549 + _T_6550; // @[Bitwise.scala 48:55:@5979.4]
  assign _T_6594 = _T_6592 + _T_6593; // @[Bitwise.scala 48:55:@5980.4]
  assign _T_6595 = _T_6591 + _T_6594; // @[Bitwise.scala 48:55:@5981.4]
  assign _T_6596 = _T_6589 + _T_6595; // @[Bitwise.scala 48:55:@5982.4]
  assign _T_6597 = _T_6584 + _T_6596; // @[Bitwise.scala 48:55:@5983.4]
  assign _T_6598 = _T_6573 + _T_6597; // @[Bitwise.scala 48:55:@5984.4]
  assign _T_6662 = _T_1124[49:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6049.4]
  assign _T_6663 = _T_6662[0]; // @[Bitwise.scala 50:65:@6050.4]
  assign _T_6664 = _T_6662[1]; // @[Bitwise.scala 50:65:@6051.4]
  assign _T_6665 = _T_6662[2]; // @[Bitwise.scala 50:65:@6052.4]
  assign _T_6666 = _T_6662[3]; // @[Bitwise.scala 50:65:@6053.4]
  assign _T_6667 = _T_6662[4]; // @[Bitwise.scala 50:65:@6054.4]
  assign _T_6668 = _T_6662[5]; // @[Bitwise.scala 50:65:@6055.4]
  assign _T_6669 = _T_6662[6]; // @[Bitwise.scala 50:65:@6056.4]
  assign _T_6670 = _T_6662[7]; // @[Bitwise.scala 50:65:@6057.4]
  assign _T_6671 = _T_6662[8]; // @[Bitwise.scala 50:65:@6058.4]
  assign _T_6672 = _T_6662[9]; // @[Bitwise.scala 50:65:@6059.4]
  assign _T_6673 = _T_6662[10]; // @[Bitwise.scala 50:65:@6060.4]
  assign _T_6674 = _T_6662[11]; // @[Bitwise.scala 50:65:@6061.4]
  assign _T_6675 = _T_6662[12]; // @[Bitwise.scala 50:65:@6062.4]
  assign _T_6676 = _T_6662[13]; // @[Bitwise.scala 50:65:@6063.4]
  assign _T_6677 = _T_6662[14]; // @[Bitwise.scala 50:65:@6064.4]
  assign _T_6678 = _T_6662[15]; // @[Bitwise.scala 50:65:@6065.4]
  assign _T_6679 = _T_6662[16]; // @[Bitwise.scala 50:65:@6066.4]
  assign _T_6680 = _T_6662[17]; // @[Bitwise.scala 50:65:@6067.4]
  assign _T_6681 = _T_6662[18]; // @[Bitwise.scala 50:65:@6068.4]
  assign _T_6682 = _T_6662[19]; // @[Bitwise.scala 50:65:@6069.4]
  assign _T_6683 = _T_6662[20]; // @[Bitwise.scala 50:65:@6070.4]
  assign _T_6684 = _T_6662[21]; // @[Bitwise.scala 50:65:@6071.4]
  assign _T_6685 = _T_6662[22]; // @[Bitwise.scala 50:65:@6072.4]
  assign _T_6686 = _T_6662[23]; // @[Bitwise.scala 50:65:@6073.4]
  assign _T_6687 = _T_6662[24]; // @[Bitwise.scala 50:65:@6074.4]
  assign _T_6688 = _T_6662[25]; // @[Bitwise.scala 50:65:@6075.4]
  assign _T_6689 = _T_6662[26]; // @[Bitwise.scala 50:65:@6076.4]
  assign _T_6690 = _T_6662[27]; // @[Bitwise.scala 50:65:@6077.4]
  assign _T_6691 = _T_6662[28]; // @[Bitwise.scala 50:65:@6078.4]
  assign _T_6692 = _T_6662[29]; // @[Bitwise.scala 50:65:@6079.4]
  assign _T_6693 = _T_6662[30]; // @[Bitwise.scala 50:65:@6080.4]
  assign _T_6694 = _T_6662[31]; // @[Bitwise.scala 50:65:@6081.4]
  assign _T_6695 = _T_6662[32]; // @[Bitwise.scala 50:65:@6082.4]
  assign _T_6696 = _T_6662[33]; // @[Bitwise.scala 50:65:@6083.4]
  assign _T_6697 = _T_6662[34]; // @[Bitwise.scala 50:65:@6084.4]
  assign _T_6698 = _T_6662[35]; // @[Bitwise.scala 50:65:@6085.4]
  assign _T_6699 = _T_6662[36]; // @[Bitwise.scala 50:65:@6086.4]
  assign _T_6700 = _T_6662[37]; // @[Bitwise.scala 50:65:@6087.4]
  assign _T_6701 = _T_6662[38]; // @[Bitwise.scala 50:65:@6088.4]
  assign _T_6702 = _T_6662[39]; // @[Bitwise.scala 50:65:@6089.4]
  assign _T_6703 = _T_6662[40]; // @[Bitwise.scala 50:65:@6090.4]
  assign _T_6704 = _T_6662[41]; // @[Bitwise.scala 50:65:@6091.4]
  assign _T_6705 = _T_6662[42]; // @[Bitwise.scala 50:65:@6092.4]
  assign _T_6706 = _T_6662[43]; // @[Bitwise.scala 50:65:@6093.4]
  assign _T_6707 = _T_6662[44]; // @[Bitwise.scala 50:65:@6094.4]
  assign _T_6708 = _T_6662[45]; // @[Bitwise.scala 50:65:@6095.4]
  assign _T_6709 = _T_6662[46]; // @[Bitwise.scala 50:65:@6096.4]
  assign _T_6710 = _T_6662[47]; // @[Bitwise.scala 50:65:@6097.4]
  assign _T_6711 = _T_6662[48]; // @[Bitwise.scala 50:65:@6098.4]
  assign _T_6712 = _T_6662[49]; // @[Bitwise.scala 50:65:@6099.4]
  assign _T_6713 = _T_6664 + _T_6665; // @[Bitwise.scala 48:55:@6100.4]
  assign _GEN_892 = {{1'd0}, _T_6663}; // @[Bitwise.scala 48:55:@6101.4]
  assign _T_6714 = _GEN_892 + _T_6713; // @[Bitwise.scala 48:55:@6101.4]
  assign _T_6715 = _T_6667 + _T_6668; // @[Bitwise.scala 48:55:@6102.4]
  assign _GEN_893 = {{1'd0}, _T_6666}; // @[Bitwise.scala 48:55:@6103.4]
  assign _T_6716 = _GEN_893 + _T_6715; // @[Bitwise.scala 48:55:@6103.4]
  assign _T_6717 = _T_6714 + _T_6716; // @[Bitwise.scala 48:55:@6104.4]
  assign _T_6718 = _T_6670 + _T_6671; // @[Bitwise.scala 48:55:@6105.4]
  assign _GEN_894 = {{1'd0}, _T_6669}; // @[Bitwise.scala 48:55:@6106.4]
  assign _T_6719 = _GEN_894 + _T_6718; // @[Bitwise.scala 48:55:@6106.4]
  assign _T_6720 = _T_6673 + _T_6674; // @[Bitwise.scala 48:55:@6107.4]
  assign _GEN_895 = {{1'd0}, _T_6672}; // @[Bitwise.scala 48:55:@6108.4]
  assign _T_6721 = _GEN_895 + _T_6720; // @[Bitwise.scala 48:55:@6108.4]
  assign _T_6722 = _T_6719 + _T_6721; // @[Bitwise.scala 48:55:@6109.4]
  assign _T_6723 = _T_6717 + _T_6722; // @[Bitwise.scala 48:55:@6110.4]
  assign _T_6724 = _T_6676 + _T_6677; // @[Bitwise.scala 48:55:@6111.4]
  assign _GEN_896 = {{1'd0}, _T_6675}; // @[Bitwise.scala 48:55:@6112.4]
  assign _T_6725 = _GEN_896 + _T_6724; // @[Bitwise.scala 48:55:@6112.4]
  assign _T_6726 = _T_6679 + _T_6680; // @[Bitwise.scala 48:55:@6113.4]
  assign _GEN_897 = {{1'd0}, _T_6678}; // @[Bitwise.scala 48:55:@6114.4]
  assign _T_6727 = _GEN_897 + _T_6726; // @[Bitwise.scala 48:55:@6114.4]
  assign _T_6728 = _T_6725 + _T_6727; // @[Bitwise.scala 48:55:@6115.4]
  assign _T_6729 = _T_6682 + _T_6683; // @[Bitwise.scala 48:55:@6116.4]
  assign _GEN_898 = {{1'd0}, _T_6681}; // @[Bitwise.scala 48:55:@6117.4]
  assign _T_6730 = _GEN_898 + _T_6729; // @[Bitwise.scala 48:55:@6117.4]
  assign _T_6731 = _T_6684 + _T_6685; // @[Bitwise.scala 48:55:@6118.4]
  assign _T_6732 = _T_6686 + _T_6687; // @[Bitwise.scala 48:55:@6119.4]
  assign _T_6733 = _T_6731 + _T_6732; // @[Bitwise.scala 48:55:@6120.4]
  assign _T_6734 = _T_6730 + _T_6733; // @[Bitwise.scala 48:55:@6121.4]
  assign _T_6735 = _T_6728 + _T_6734; // @[Bitwise.scala 48:55:@6122.4]
  assign _T_6736 = _T_6723 + _T_6735; // @[Bitwise.scala 48:55:@6123.4]
  assign _T_6737 = _T_6689 + _T_6690; // @[Bitwise.scala 48:55:@6124.4]
  assign _GEN_899 = {{1'd0}, _T_6688}; // @[Bitwise.scala 48:55:@6125.4]
  assign _T_6738 = _GEN_899 + _T_6737; // @[Bitwise.scala 48:55:@6125.4]
  assign _T_6739 = _T_6692 + _T_6693; // @[Bitwise.scala 48:55:@6126.4]
  assign _GEN_900 = {{1'd0}, _T_6691}; // @[Bitwise.scala 48:55:@6127.4]
  assign _T_6740 = _GEN_900 + _T_6739; // @[Bitwise.scala 48:55:@6127.4]
  assign _T_6741 = _T_6738 + _T_6740; // @[Bitwise.scala 48:55:@6128.4]
  assign _T_6742 = _T_6695 + _T_6696; // @[Bitwise.scala 48:55:@6129.4]
  assign _GEN_901 = {{1'd0}, _T_6694}; // @[Bitwise.scala 48:55:@6130.4]
  assign _T_6743 = _GEN_901 + _T_6742; // @[Bitwise.scala 48:55:@6130.4]
  assign _T_6744 = _T_6698 + _T_6699; // @[Bitwise.scala 48:55:@6131.4]
  assign _GEN_902 = {{1'd0}, _T_6697}; // @[Bitwise.scala 48:55:@6132.4]
  assign _T_6745 = _GEN_902 + _T_6744; // @[Bitwise.scala 48:55:@6132.4]
  assign _T_6746 = _T_6743 + _T_6745; // @[Bitwise.scala 48:55:@6133.4]
  assign _T_6747 = _T_6741 + _T_6746; // @[Bitwise.scala 48:55:@6134.4]
  assign _T_6748 = _T_6701 + _T_6702; // @[Bitwise.scala 48:55:@6135.4]
  assign _GEN_903 = {{1'd0}, _T_6700}; // @[Bitwise.scala 48:55:@6136.4]
  assign _T_6749 = _GEN_903 + _T_6748; // @[Bitwise.scala 48:55:@6136.4]
  assign _T_6750 = _T_6704 + _T_6705; // @[Bitwise.scala 48:55:@6137.4]
  assign _GEN_904 = {{1'd0}, _T_6703}; // @[Bitwise.scala 48:55:@6138.4]
  assign _T_6751 = _GEN_904 + _T_6750; // @[Bitwise.scala 48:55:@6138.4]
  assign _T_6752 = _T_6749 + _T_6751; // @[Bitwise.scala 48:55:@6139.4]
  assign _T_6753 = _T_6707 + _T_6708; // @[Bitwise.scala 48:55:@6140.4]
  assign _GEN_905 = {{1'd0}, _T_6706}; // @[Bitwise.scala 48:55:@6141.4]
  assign _T_6754 = _GEN_905 + _T_6753; // @[Bitwise.scala 48:55:@6141.4]
  assign _T_6755 = _T_6709 + _T_6710; // @[Bitwise.scala 48:55:@6142.4]
  assign _T_6756 = _T_6711 + _T_6712; // @[Bitwise.scala 48:55:@6143.4]
  assign _T_6757 = _T_6755 + _T_6756; // @[Bitwise.scala 48:55:@6144.4]
  assign _T_6758 = _T_6754 + _T_6757; // @[Bitwise.scala 48:55:@6145.4]
  assign _T_6759 = _T_6752 + _T_6758; // @[Bitwise.scala 48:55:@6146.4]
  assign _T_6760 = _T_6747 + _T_6759; // @[Bitwise.scala 48:55:@6147.4]
  assign _T_6761 = _T_6736 + _T_6760; // @[Bitwise.scala 48:55:@6148.4]
  assign _T_6825 = _T_1124[50:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6213.4]
  assign _T_6826 = _T_6825[0]; // @[Bitwise.scala 50:65:@6214.4]
  assign _T_6827 = _T_6825[1]; // @[Bitwise.scala 50:65:@6215.4]
  assign _T_6828 = _T_6825[2]; // @[Bitwise.scala 50:65:@6216.4]
  assign _T_6829 = _T_6825[3]; // @[Bitwise.scala 50:65:@6217.4]
  assign _T_6830 = _T_6825[4]; // @[Bitwise.scala 50:65:@6218.4]
  assign _T_6831 = _T_6825[5]; // @[Bitwise.scala 50:65:@6219.4]
  assign _T_6832 = _T_6825[6]; // @[Bitwise.scala 50:65:@6220.4]
  assign _T_6833 = _T_6825[7]; // @[Bitwise.scala 50:65:@6221.4]
  assign _T_6834 = _T_6825[8]; // @[Bitwise.scala 50:65:@6222.4]
  assign _T_6835 = _T_6825[9]; // @[Bitwise.scala 50:65:@6223.4]
  assign _T_6836 = _T_6825[10]; // @[Bitwise.scala 50:65:@6224.4]
  assign _T_6837 = _T_6825[11]; // @[Bitwise.scala 50:65:@6225.4]
  assign _T_6838 = _T_6825[12]; // @[Bitwise.scala 50:65:@6226.4]
  assign _T_6839 = _T_6825[13]; // @[Bitwise.scala 50:65:@6227.4]
  assign _T_6840 = _T_6825[14]; // @[Bitwise.scala 50:65:@6228.4]
  assign _T_6841 = _T_6825[15]; // @[Bitwise.scala 50:65:@6229.4]
  assign _T_6842 = _T_6825[16]; // @[Bitwise.scala 50:65:@6230.4]
  assign _T_6843 = _T_6825[17]; // @[Bitwise.scala 50:65:@6231.4]
  assign _T_6844 = _T_6825[18]; // @[Bitwise.scala 50:65:@6232.4]
  assign _T_6845 = _T_6825[19]; // @[Bitwise.scala 50:65:@6233.4]
  assign _T_6846 = _T_6825[20]; // @[Bitwise.scala 50:65:@6234.4]
  assign _T_6847 = _T_6825[21]; // @[Bitwise.scala 50:65:@6235.4]
  assign _T_6848 = _T_6825[22]; // @[Bitwise.scala 50:65:@6236.4]
  assign _T_6849 = _T_6825[23]; // @[Bitwise.scala 50:65:@6237.4]
  assign _T_6850 = _T_6825[24]; // @[Bitwise.scala 50:65:@6238.4]
  assign _T_6851 = _T_6825[25]; // @[Bitwise.scala 50:65:@6239.4]
  assign _T_6852 = _T_6825[26]; // @[Bitwise.scala 50:65:@6240.4]
  assign _T_6853 = _T_6825[27]; // @[Bitwise.scala 50:65:@6241.4]
  assign _T_6854 = _T_6825[28]; // @[Bitwise.scala 50:65:@6242.4]
  assign _T_6855 = _T_6825[29]; // @[Bitwise.scala 50:65:@6243.4]
  assign _T_6856 = _T_6825[30]; // @[Bitwise.scala 50:65:@6244.4]
  assign _T_6857 = _T_6825[31]; // @[Bitwise.scala 50:65:@6245.4]
  assign _T_6858 = _T_6825[32]; // @[Bitwise.scala 50:65:@6246.4]
  assign _T_6859 = _T_6825[33]; // @[Bitwise.scala 50:65:@6247.4]
  assign _T_6860 = _T_6825[34]; // @[Bitwise.scala 50:65:@6248.4]
  assign _T_6861 = _T_6825[35]; // @[Bitwise.scala 50:65:@6249.4]
  assign _T_6862 = _T_6825[36]; // @[Bitwise.scala 50:65:@6250.4]
  assign _T_6863 = _T_6825[37]; // @[Bitwise.scala 50:65:@6251.4]
  assign _T_6864 = _T_6825[38]; // @[Bitwise.scala 50:65:@6252.4]
  assign _T_6865 = _T_6825[39]; // @[Bitwise.scala 50:65:@6253.4]
  assign _T_6866 = _T_6825[40]; // @[Bitwise.scala 50:65:@6254.4]
  assign _T_6867 = _T_6825[41]; // @[Bitwise.scala 50:65:@6255.4]
  assign _T_6868 = _T_6825[42]; // @[Bitwise.scala 50:65:@6256.4]
  assign _T_6869 = _T_6825[43]; // @[Bitwise.scala 50:65:@6257.4]
  assign _T_6870 = _T_6825[44]; // @[Bitwise.scala 50:65:@6258.4]
  assign _T_6871 = _T_6825[45]; // @[Bitwise.scala 50:65:@6259.4]
  assign _T_6872 = _T_6825[46]; // @[Bitwise.scala 50:65:@6260.4]
  assign _T_6873 = _T_6825[47]; // @[Bitwise.scala 50:65:@6261.4]
  assign _T_6874 = _T_6825[48]; // @[Bitwise.scala 50:65:@6262.4]
  assign _T_6875 = _T_6825[49]; // @[Bitwise.scala 50:65:@6263.4]
  assign _T_6876 = _T_6825[50]; // @[Bitwise.scala 50:65:@6264.4]
  assign _T_6877 = _T_6827 + _T_6828; // @[Bitwise.scala 48:55:@6265.4]
  assign _GEN_906 = {{1'd0}, _T_6826}; // @[Bitwise.scala 48:55:@6266.4]
  assign _T_6878 = _GEN_906 + _T_6877; // @[Bitwise.scala 48:55:@6266.4]
  assign _T_6879 = _T_6830 + _T_6831; // @[Bitwise.scala 48:55:@6267.4]
  assign _GEN_907 = {{1'd0}, _T_6829}; // @[Bitwise.scala 48:55:@6268.4]
  assign _T_6880 = _GEN_907 + _T_6879; // @[Bitwise.scala 48:55:@6268.4]
  assign _T_6881 = _T_6878 + _T_6880; // @[Bitwise.scala 48:55:@6269.4]
  assign _T_6882 = _T_6833 + _T_6834; // @[Bitwise.scala 48:55:@6270.4]
  assign _GEN_908 = {{1'd0}, _T_6832}; // @[Bitwise.scala 48:55:@6271.4]
  assign _T_6883 = _GEN_908 + _T_6882; // @[Bitwise.scala 48:55:@6271.4]
  assign _T_6884 = _T_6836 + _T_6837; // @[Bitwise.scala 48:55:@6272.4]
  assign _GEN_909 = {{1'd0}, _T_6835}; // @[Bitwise.scala 48:55:@6273.4]
  assign _T_6885 = _GEN_909 + _T_6884; // @[Bitwise.scala 48:55:@6273.4]
  assign _T_6886 = _T_6883 + _T_6885; // @[Bitwise.scala 48:55:@6274.4]
  assign _T_6887 = _T_6881 + _T_6886; // @[Bitwise.scala 48:55:@6275.4]
  assign _T_6888 = _T_6839 + _T_6840; // @[Bitwise.scala 48:55:@6276.4]
  assign _GEN_910 = {{1'd0}, _T_6838}; // @[Bitwise.scala 48:55:@6277.4]
  assign _T_6889 = _GEN_910 + _T_6888; // @[Bitwise.scala 48:55:@6277.4]
  assign _T_6890 = _T_6842 + _T_6843; // @[Bitwise.scala 48:55:@6278.4]
  assign _GEN_911 = {{1'd0}, _T_6841}; // @[Bitwise.scala 48:55:@6279.4]
  assign _T_6891 = _GEN_911 + _T_6890; // @[Bitwise.scala 48:55:@6279.4]
  assign _T_6892 = _T_6889 + _T_6891; // @[Bitwise.scala 48:55:@6280.4]
  assign _T_6893 = _T_6845 + _T_6846; // @[Bitwise.scala 48:55:@6281.4]
  assign _GEN_912 = {{1'd0}, _T_6844}; // @[Bitwise.scala 48:55:@6282.4]
  assign _T_6894 = _GEN_912 + _T_6893; // @[Bitwise.scala 48:55:@6282.4]
  assign _T_6895 = _T_6847 + _T_6848; // @[Bitwise.scala 48:55:@6283.4]
  assign _T_6896 = _T_6849 + _T_6850; // @[Bitwise.scala 48:55:@6284.4]
  assign _T_6897 = _T_6895 + _T_6896; // @[Bitwise.scala 48:55:@6285.4]
  assign _T_6898 = _T_6894 + _T_6897; // @[Bitwise.scala 48:55:@6286.4]
  assign _T_6899 = _T_6892 + _T_6898; // @[Bitwise.scala 48:55:@6287.4]
  assign _T_6900 = _T_6887 + _T_6899; // @[Bitwise.scala 48:55:@6288.4]
  assign _T_6901 = _T_6852 + _T_6853; // @[Bitwise.scala 48:55:@6289.4]
  assign _GEN_913 = {{1'd0}, _T_6851}; // @[Bitwise.scala 48:55:@6290.4]
  assign _T_6902 = _GEN_913 + _T_6901; // @[Bitwise.scala 48:55:@6290.4]
  assign _T_6903 = _T_6855 + _T_6856; // @[Bitwise.scala 48:55:@6291.4]
  assign _GEN_914 = {{1'd0}, _T_6854}; // @[Bitwise.scala 48:55:@6292.4]
  assign _T_6904 = _GEN_914 + _T_6903; // @[Bitwise.scala 48:55:@6292.4]
  assign _T_6905 = _T_6902 + _T_6904; // @[Bitwise.scala 48:55:@6293.4]
  assign _T_6906 = _T_6858 + _T_6859; // @[Bitwise.scala 48:55:@6294.4]
  assign _GEN_915 = {{1'd0}, _T_6857}; // @[Bitwise.scala 48:55:@6295.4]
  assign _T_6907 = _GEN_915 + _T_6906; // @[Bitwise.scala 48:55:@6295.4]
  assign _T_6908 = _T_6860 + _T_6861; // @[Bitwise.scala 48:55:@6296.4]
  assign _T_6909 = _T_6862 + _T_6863; // @[Bitwise.scala 48:55:@6297.4]
  assign _T_6910 = _T_6908 + _T_6909; // @[Bitwise.scala 48:55:@6298.4]
  assign _T_6911 = _T_6907 + _T_6910; // @[Bitwise.scala 48:55:@6299.4]
  assign _T_6912 = _T_6905 + _T_6911; // @[Bitwise.scala 48:55:@6300.4]
  assign _T_6913 = _T_6865 + _T_6866; // @[Bitwise.scala 48:55:@6301.4]
  assign _GEN_916 = {{1'd0}, _T_6864}; // @[Bitwise.scala 48:55:@6302.4]
  assign _T_6914 = _GEN_916 + _T_6913; // @[Bitwise.scala 48:55:@6302.4]
  assign _T_6915 = _T_6868 + _T_6869; // @[Bitwise.scala 48:55:@6303.4]
  assign _GEN_917 = {{1'd0}, _T_6867}; // @[Bitwise.scala 48:55:@6304.4]
  assign _T_6916 = _GEN_917 + _T_6915; // @[Bitwise.scala 48:55:@6304.4]
  assign _T_6917 = _T_6914 + _T_6916; // @[Bitwise.scala 48:55:@6305.4]
  assign _T_6918 = _T_6871 + _T_6872; // @[Bitwise.scala 48:55:@6306.4]
  assign _GEN_918 = {{1'd0}, _T_6870}; // @[Bitwise.scala 48:55:@6307.4]
  assign _T_6919 = _GEN_918 + _T_6918; // @[Bitwise.scala 48:55:@6307.4]
  assign _T_6920 = _T_6873 + _T_6874; // @[Bitwise.scala 48:55:@6308.4]
  assign _T_6921 = _T_6875 + _T_6876; // @[Bitwise.scala 48:55:@6309.4]
  assign _T_6922 = _T_6920 + _T_6921; // @[Bitwise.scala 48:55:@6310.4]
  assign _T_6923 = _T_6919 + _T_6922; // @[Bitwise.scala 48:55:@6311.4]
  assign _T_6924 = _T_6917 + _T_6923; // @[Bitwise.scala 48:55:@6312.4]
  assign _T_6925 = _T_6912 + _T_6924; // @[Bitwise.scala 48:55:@6313.4]
  assign _T_6926 = _T_6900 + _T_6925; // @[Bitwise.scala 48:55:@6314.4]
  assign _T_6990 = _T_1124[51:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6379.4]
  assign _T_6991 = _T_6990[0]; // @[Bitwise.scala 50:65:@6380.4]
  assign _T_6992 = _T_6990[1]; // @[Bitwise.scala 50:65:@6381.4]
  assign _T_6993 = _T_6990[2]; // @[Bitwise.scala 50:65:@6382.4]
  assign _T_6994 = _T_6990[3]; // @[Bitwise.scala 50:65:@6383.4]
  assign _T_6995 = _T_6990[4]; // @[Bitwise.scala 50:65:@6384.4]
  assign _T_6996 = _T_6990[5]; // @[Bitwise.scala 50:65:@6385.4]
  assign _T_6997 = _T_6990[6]; // @[Bitwise.scala 50:65:@6386.4]
  assign _T_6998 = _T_6990[7]; // @[Bitwise.scala 50:65:@6387.4]
  assign _T_6999 = _T_6990[8]; // @[Bitwise.scala 50:65:@6388.4]
  assign _T_7000 = _T_6990[9]; // @[Bitwise.scala 50:65:@6389.4]
  assign _T_7001 = _T_6990[10]; // @[Bitwise.scala 50:65:@6390.4]
  assign _T_7002 = _T_6990[11]; // @[Bitwise.scala 50:65:@6391.4]
  assign _T_7003 = _T_6990[12]; // @[Bitwise.scala 50:65:@6392.4]
  assign _T_7004 = _T_6990[13]; // @[Bitwise.scala 50:65:@6393.4]
  assign _T_7005 = _T_6990[14]; // @[Bitwise.scala 50:65:@6394.4]
  assign _T_7006 = _T_6990[15]; // @[Bitwise.scala 50:65:@6395.4]
  assign _T_7007 = _T_6990[16]; // @[Bitwise.scala 50:65:@6396.4]
  assign _T_7008 = _T_6990[17]; // @[Bitwise.scala 50:65:@6397.4]
  assign _T_7009 = _T_6990[18]; // @[Bitwise.scala 50:65:@6398.4]
  assign _T_7010 = _T_6990[19]; // @[Bitwise.scala 50:65:@6399.4]
  assign _T_7011 = _T_6990[20]; // @[Bitwise.scala 50:65:@6400.4]
  assign _T_7012 = _T_6990[21]; // @[Bitwise.scala 50:65:@6401.4]
  assign _T_7013 = _T_6990[22]; // @[Bitwise.scala 50:65:@6402.4]
  assign _T_7014 = _T_6990[23]; // @[Bitwise.scala 50:65:@6403.4]
  assign _T_7015 = _T_6990[24]; // @[Bitwise.scala 50:65:@6404.4]
  assign _T_7016 = _T_6990[25]; // @[Bitwise.scala 50:65:@6405.4]
  assign _T_7017 = _T_6990[26]; // @[Bitwise.scala 50:65:@6406.4]
  assign _T_7018 = _T_6990[27]; // @[Bitwise.scala 50:65:@6407.4]
  assign _T_7019 = _T_6990[28]; // @[Bitwise.scala 50:65:@6408.4]
  assign _T_7020 = _T_6990[29]; // @[Bitwise.scala 50:65:@6409.4]
  assign _T_7021 = _T_6990[30]; // @[Bitwise.scala 50:65:@6410.4]
  assign _T_7022 = _T_6990[31]; // @[Bitwise.scala 50:65:@6411.4]
  assign _T_7023 = _T_6990[32]; // @[Bitwise.scala 50:65:@6412.4]
  assign _T_7024 = _T_6990[33]; // @[Bitwise.scala 50:65:@6413.4]
  assign _T_7025 = _T_6990[34]; // @[Bitwise.scala 50:65:@6414.4]
  assign _T_7026 = _T_6990[35]; // @[Bitwise.scala 50:65:@6415.4]
  assign _T_7027 = _T_6990[36]; // @[Bitwise.scala 50:65:@6416.4]
  assign _T_7028 = _T_6990[37]; // @[Bitwise.scala 50:65:@6417.4]
  assign _T_7029 = _T_6990[38]; // @[Bitwise.scala 50:65:@6418.4]
  assign _T_7030 = _T_6990[39]; // @[Bitwise.scala 50:65:@6419.4]
  assign _T_7031 = _T_6990[40]; // @[Bitwise.scala 50:65:@6420.4]
  assign _T_7032 = _T_6990[41]; // @[Bitwise.scala 50:65:@6421.4]
  assign _T_7033 = _T_6990[42]; // @[Bitwise.scala 50:65:@6422.4]
  assign _T_7034 = _T_6990[43]; // @[Bitwise.scala 50:65:@6423.4]
  assign _T_7035 = _T_6990[44]; // @[Bitwise.scala 50:65:@6424.4]
  assign _T_7036 = _T_6990[45]; // @[Bitwise.scala 50:65:@6425.4]
  assign _T_7037 = _T_6990[46]; // @[Bitwise.scala 50:65:@6426.4]
  assign _T_7038 = _T_6990[47]; // @[Bitwise.scala 50:65:@6427.4]
  assign _T_7039 = _T_6990[48]; // @[Bitwise.scala 50:65:@6428.4]
  assign _T_7040 = _T_6990[49]; // @[Bitwise.scala 50:65:@6429.4]
  assign _T_7041 = _T_6990[50]; // @[Bitwise.scala 50:65:@6430.4]
  assign _T_7042 = _T_6990[51]; // @[Bitwise.scala 50:65:@6431.4]
  assign _T_7043 = _T_6992 + _T_6993; // @[Bitwise.scala 48:55:@6432.4]
  assign _GEN_919 = {{1'd0}, _T_6991}; // @[Bitwise.scala 48:55:@6433.4]
  assign _T_7044 = _GEN_919 + _T_7043; // @[Bitwise.scala 48:55:@6433.4]
  assign _T_7045 = _T_6995 + _T_6996; // @[Bitwise.scala 48:55:@6434.4]
  assign _GEN_920 = {{1'd0}, _T_6994}; // @[Bitwise.scala 48:55:@6435.4]
  assign _T_7046 = _GEN_920 + _T_7045; // @[Bitwise.scala 48:55:@6435.4]
  assign _T_7047 = _T_7044 + _T_7046; // @[Bitwise.scala 48:55:@6436.4]
  assign _T_7048 = _T_6998 + _T_6999; // @[Bitwise.scala 48:55:@6437.4]
  assign _GEN_921 = {{1'd0}, _T_6997}; // @[Bitwise.scala 48:55:@6438.4]
  assign _T_7049 = _GEN_921 + _T_7048; // @[Bitwise.scala 48:55:@6438.4]
  assign _T_7050 = _T_7000 + _T_7001; // @[Bitwise.scala 48:55:@6439.4]
  assign _T_7051 = _T_7002 + _T_7003; // @[Bitwise.scala 48:55:@6440.4]
  assign _T_7052 = _T_7050 + _T_7051; // @[Bitwise.scala 48:55:@6441.4]
  assign _T_7053 = _T_7049 + _T_7052; // @[Bitwise.scala 48:55:@6442.4]
  assign _T_7054 = _T_7047 + _T_7053; // @[Bitwise.scala 48:55:@6443.4]
  assign _T_7055 = _T_7005 + _T_7006; // @[Bitwise.scala 48:55:@6444.4]
  assign _GEN_922 = {{1'd0}, _T_7004}; // @[Bitwise.scala 48:55:@6445.4]
  assign _T_7056 = _GEN_922 + _T_7055; // @[Bitwise.scala 48:55:@6445.4]
  assign _T_7057 = _T_7008 + _T_7009; // @[Bitwise.scala 48:55:@6446.4]
  assign _GEN_923 = {{1'd0}, _T_7007}; // @[Bitwise.scala 48:55:@6447.4]
  assign _T_7058 = _GEN_923 + _T_7057; // @[Bitwise.scala 48:55:@6447.4]
  assign _T_7059 = _T_7056 + _T_7058; // @[Bitwise.scala 48:55:@6448.4]
  assign _T_7060 = _T_7011 + _T_7012; // @[Bitwise.scala 48:55:@6449.4]
  assign _GEN_924 = {{1'd0}, _T_7010}; // @[Bitwise.scala 48:55:@6450.4]
  assign _T_7061 = _GEN_924 + _T_7060; // @[Bitwise.scala 48:55:@6450.4]
  assign _T_7062 = _T_7013 + _T_7014; // @[Bitwise.scala 48:55:@6451.4]
  assign _T_7063 = _T_7015 + _T_7016; // @[Bitwise.scala 48:55:@6452.4]
  assign _T_7064 = _T_7062 + _T_7063; // @[Bitwise.scala 48:55:@6453.4]
  assign _T_7065 = _T_7061 + _T_7064; // @[Bitwise.scala 48:55:@6454.4]
  assign _T_7066 = _T_7059 + _T_7065; // @[Bitwise.scala 48:55:@6455.4]
  assign _T_7067 = _T_7054 + _T_7066; // @[Bitwise.scala 48:55:@6456.4]
  assign _T_7068 = _T_7018 + _T_7019; // @[Bitwise.scala 48:55:@6457.4]
  assign _GEN_925 = {{1'd0}, _T_7017}; // @[Bitwise.scala 48:55:@6458.4]
  assign _T_7069 = _GEN_925 + _T_7068; // @[Bitwise.scala 48:55:@6458.4]
  assign _T_7070 = _T_7021 + _T_7022; // @[Bitwise.scala 48:55:@6459.4]
  assign _GEN_926 = {{1'd0}, _T_7020}; // @[Bitwise.scala 48:55:@6460.4]
  assign _T_7071 = _GEN_926 + _T_7070; // @[Bitwise.scala 48:55:@6460.4]
  assign _T_7072 = _T_7069 + _T_7071; // @[Bitwise.scala 48:55:@6461.4]
  assign _T_7073 = _T_7024 + _T_7025; // @[Bitwise.scala 48:55:@6462.4]
  assign _GEN_927 = {{1'd0}, _T_7023}; // @[Bitwise.scala 48:55:@6463.4]
  assign _T_7074 = _GEN_927 + _T_7073; // @[Bitwise.scala 48:55:@6463.4]
  assign _T_7075 = _T_7026 + _T_7027; // @[Bitwise.scala 48:55:@6464.4]
  assign _T_7076 = _T_7028 + _T_7029; // @[Bitwise.scala 48:55:@6465.4]
  assign _T_7077 = _T_7075 + _T_7076; // @[Bitwise.scala 48:55:@6466.4]
  assign _T_7078 = _T_7074 + _T_7077; // @[Bitwise.scala 48:55:@6467.4]
  assign _T_7079 = _T_7072 + _T_7078; // @[Bitwise.scala 48:55:@6468.4]
  assign _T_7080 = _T_7031 + _T_7032; // @[Bitwise.scala 48:55:@6469.4]
  assign _GEN_928 = {{1'd0}, _T_7030}; // @[Bitwise.scala 48:55:@6470.4]
  assign _T_7081 = _GEN_928 + _T_7080; // @[Bitwise.scala 48:55:@6470.4]
  assign _T_7082 = _T_7034 + _T_7035; // @[Bitwise.scala 48:55:@6471.4]
  assign _GEN_929 = {{1'd0}, _T_7033}; // @[Bitwise.scala 48:55:@6472.4]
  assign _T_7083 = _GEN_929 + _T_7082; // @[Bitwise.scala 48:55:@6472.4]
  assign _T_7084 = _T_7081 + _T_7083; // @[Bitwise.scala 48:55:@6473.4]
  assign _T_7085 = _T_7037 + _T_7038; // @[Bitwise.scala 48:55:@6474.4]
  assign _GEN_930 = {{1'd0}, _T_7036}; // @[Bitwise.scala 48:55:@6475.4]
  assign _T_7086 = _GEN_930 + _T_7085; // @[Bitwise.scala 48:55:@6475.4]
  assign _T_7087 = _T_7039 + _T_7040; // @[Bitwise.scala 48:55:@6476.4]
  assign _T_7088 = _T_7041 + _T_7042; // @[Bitwise.scala 48:55:@6477.4]
  assign _T_7089 = _T_7087 + _T_7088; // @[Bitwise.scala 48:55:@6478.4]
  assign _T_7090 = _T_7086 + _T_7089; // @[Bitwise.scala 48:55:@6479.4]
  assign _T_7091 = _T_7084 + _T_7090; // @[Bitwise.scala 48:55:@6480.4]
  assign _T_7092 = _T_7079 + _T_7091; // @[Bitwise.scala 48:55:@6481.4]
  assign _T_7093 = _T_7067 + _T_7092; // @[Bitwise.scala 48:55:@6482.4]
  assign _T_7157 = _T_1124[52:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6547.4]
  assign _T_7158 = _T_7157[0]; // @[Bitwise.scala 50:65:@6548.4]
  assign _T_7159 = _T_7157[1]; // @[Bitwise.scala 50:65:@6549.4]
  assign _T_7160 = _T_7157[2]; // @[Bitwise.scala 50:65:@6550.4]
  assign _T_7161 = _T_7157[3]; // @[Bitwise.scala 50:65:@6551.4]
  assign _T_7162 = _T_7157[4]; // @[Bitwise.scala 50:65:@6552.4]
  assign _T_7163 = _T_7157[5]; // @[Bitwise.scala 50:65:@6553.4]
  assign _T_7164 = _T_7157[6]; // @[Bitwise.scala 50:65:@6554.4]
  assign _T_7165 = _T_7157[7]; // @[Bitwise.scala 50:65:@6555.4]
  assign _T_7166 = _T_7157[8]; // @[Bitwise.scala 50:65:@6556.4]
  assign _T_7167 = _T_7157[9]; // @[Bitwise.scala 50:65:@6557.4]
  assign _T_7168 = _T_7157[10]; // @[Bitwise.scala 50:65:@6558.4]
  assign _T_7169 = _T_7157[11]; // @[Bitwise.scala 50:65:@6559.4]
  assign _T_7170 = _T_7157[12]; // @[Bitwise.scala 50:65:@6560.4]
  assign _T_7171 = _T_7157[13]; // @[Bitwise.scala 50:65:@6561.4]
  assign _T_7172 = _T_7157[14]; // @[Bitwise.scala 50:65:@6562.4]
  assign _T_7173 = _T_7157[15]; // @[Bitwise.scala 50:65:@6563.4]
  assign _T_7174 = _T_7157[16]; // @[Bitwise.scala 50:65:@6564.4]
  assign _T_7175 = _T_7157[17]; // @[Bitwise.scala 50:65:@6565.4]
  assign _T_7176 = _T_7157[18]; // @[Bitwise.scala 50:65:@6566.4]
  assign _T_7177 = _T_7157[19]; // @[Bitwise.scala 50:65:@6567.4]
  assign _T_7178 = _T_7157[20]; // @[Bitwise.scala 50:65:@6568.4]
  assign _T_7179 = _T_7157[21]; // @[Bitwise.scala 50:65:@6569.4]
  assign _T_7180 = _T_7157[22]; // @[Bitwise.scala 50:65:@6570.4]
  assign _T_7181 = _T_7157[23]; // @[Bitwise.scala 50:65:@6571.4]
  assign _T_7182 = _T_7157[24]; // @[Bitwise.scala 50:65:@6572.4]
  assign _T_7183 = _T_7157[25]; // @[Bitwise.scala 50:65:@6573.4]
  assign _T_7184 = _T_7157[26]; // @[Bitwise.scala 50:65:@6574.4]
  assign _T_7185 = _T_7157[27]; // @[Bitwise.scala 50:65:@6575.4]
  assign _T_7186 = _T_7157[28]; // @[Bitwise.scala 50:65:@6576.4]
  assign _T_7187 = _T_7157[29]; // @[Bitwise.scala 50:65:@6577.4]
  assign _T_7188 = _T_7157[30]; // @[Bitwise.scala 50:65:@6578.4]
  assign _T_7189 = _T_7157[31]; // @[Bitwise.scala 50:65:@6579.4]
  assign _T_7190 = _T_7157[32]; // @[Bitwise.scala 50:65:@6580.4]
  assign _T_7191 = _T_7157[33]; // @[Bitwise.scala 50:65:@6581.4]
  assign _T_7192 = _T_7157[34]; // @[Bitwise.scala 50:65:@6582.4]
  assign _T_7193 = _T_7157[35]; // @[Bitwise.scala 50:65:@6583.4]
  assign _T_7194 = _T_7157[36]; // @[Bitwise.scala 50:65:@6584.4]
  assign _T_7195 = _T_7157[37]; // @[Bitwise.scala 50:65:@6585.4]
  assign _T_7196 = _T_7157[38]; // @[Bitwise.scala 50:65:@6586.4]
  assign _T_7197 = _T_7157[39]; // @[Bitwise.scala 50:65:@6587.4]
  assign _T_7198 = _T_7157[40]; // @[Bitwise.scala 50:65:@6588.4]
  assign _T_7199 = _T_7157[41]; // @[Bitwise.scala 50:65:@6589.4]
  assign _T_7200 = _T_7157[42]; // @[Bitwise.scala 50:65:@6590.4]
  assign _T_7201 = _T_7157[43]; // @[Bitwise.scala 50:65:@6591.4]
  assign _T_7202 = _T_7157[44]; // @[Bitwise.scala 50:65:@6592.4]
  assign _T_7203 = _T_7157[45]; // @[Bitwise.scala 50:65:@6593.4]
  assign _T_7204 = _T_7157[46]; // @[Bitwise.scala 50:65:@6594.4]
  assign _T_7205 = _T_7157[47]; // @[Bitwise.scala 50:65:@6595.4]
  assign _T_7206 = _T_7157[48]; // @[Bitwise.scala 50:65:@6596.4]
  assign _T_7207 = _T_7157[49]; // @[Bitwise.scala 50:65:@6597.4]
  assign _T_7208 = _T_7157[50]; // @[Bitwise.scala 50:65:@6598.4]
  assign _T_7209 = _T_7157[51]; // @[Bitwise.scala 50:65:@6599.4]
  assign _T_7210 = _T_7157[52]; // @[Bitwise.scala 50:65:@6600.4]
  assign _T_7211 = _T_7159 + _T_7160; // @[Bitwise.scala 48:55:@6601.4]
  assign _GEN_931 = {{1'd0}, _T_7158}; // @[Bitwise.scala 48:55:@6602.4]
  assign _T_7212 = _GEN_931 + _T_7211; // @[Bitwise.scala 48:55:@6602.4]
  assign _T_7213 = _T_7162 + _T_7163; // @[Bitwise.scala 48:55:@6603.4]
  assign _GEN_932 = {{1'd0}, _T_7161}; // @[Bitwise.scala 48:55:@6604.4]
  assign _T_7214 = _GEN_932 + _T_7213; // @[Bitwise.scala 48:55:@6604.4]
  assign _T_7215 = _T_7212 + _T_7214; // @[Bitwise.scala 48:55:@6605.4]
  assign _T_7216 = _T_7165 + _T_7166; // @[Bitwise.scala 48:55:@6606.4]
  assign _GEN_933 = {{1'd0}, _T_7164}; // @[Bitwise.scala 48:55:@6607.4]
  assign _T_7217 = _GEN_933 + _T_7216; // @[Bitwise.scala 48:55:@6607.4]
  assign _T_7218 = _T_7167 + _T_7168; // @[Bitwise.scala 48:55:@6608.4]
  assign _T_7219 = _T_7169 + _T_7170; // @[Bitwise.scala 48:55:@6609.4]
  assign _T_7220 = _T_7218 + _T_7219; // @[Bitwise.scala 48:55:@6610.4]
  assign _T_7221 = _T_7217 + _T_7220; // @[Bitwise.scala 48:55:@6611.4]
  assign _T_7222 = _T_7215 + _T_7221; // @[Bitwise.scala 48:55:@6612.4]
  assign _T_7223 = _T_7172 + _T_7173; // @[Bitwise.scala 48:55:@6613.4]
  assign _GEN_934 = {{1'd0}, _T_7171}; // @[Bitwise.scala 48:55:@6614.4]
  assign _T_7224 = _GEN_934 + _T_7223; // @[Bitwise.scala 48:55:@6614.4]
  assign _T_7225 = _T_7175 + _T_7176; // @[Bitwise.scala 48:55:@6615.4]
  assign _GEN_935 = {{1'd0}, _T_7174}; // @[Bitwise.scala 48:55:@6616.4]
  assign _T_7226 = _GEN_935 + _T_7225; // @[Bitwise.scala 48:55:@6616.4]
  assign _T_7227 = _T_7224 + _T_7226; // @[Bitwise.scala 48:55:@6617.4]
  assign _T_7228 = _T_7178 + _T_7179; // @[Bitwise.scala 48:55:@6618.4]
  assign _GEN_936 = {{1'd0}, _T_7177}; // @[Bitwise.scala 48:55:@6619.4]
  assign _T_7229 = _GEN_936 + _T_7228; // @[Bitwise.scala 48:55:@6619.4]
  assign _T_7230 = _T_7180 + _T_7181; // @[Bitwise.scala 48:55:@6620.4]
  assign _T_7231 = _T_7182 + _T_7183; // @[Bitwise.scala 48:55:@6621.4]
  assign _T_7232 = _T_7230 + _T_7231; // @[Bitwise.scala 48:55:@6622.4]
  assign _T_7233 = _T_7229 + _T_7232; // @[Bitwise.scala 48:55:@6623.4]
  assign _T_7234 = _T_7227 + _T_7233; // @[Bitwise.scala 48:55:@6624.4]
  assign _T_7235 = _T_7222 + _T_7234; // @[Bitwise.scala 48:55:@6625.4]
  assign _T_7236 = _T_7185 + _T_7186; // @[Bitwise.scala 48:55:@6626.4]
  assign _GEN_937 = {{1'd0}, _T_7184}; // @[Bitwise.scala 48:55:@6627.4]
  assign _T_7237 = _GEN_937 + _T_7236; // @[Bitwise.scala 48:55:@6627.4]
  assign _T_7238 = _T_7188 + _T_7189; // @[Bitwise.scala 48:55:@6628.4]
  assign _GEN_938 = {{1'd0}, _T_7187}; // @[Bitwise.scala 48:55:@6629.4]
  assign _T_7239 = _GEN_938 + _T_7238; // @[Bitwise.scala 48:55:@6629.4]
  assign _T_7240 = _T_7237 + _T_7239; // @[Bitwise.scala 48:55:@6630.4]
  assign _T_7241 = _T_7191 + _T_7192; // @[Bitwise.scala 48:55:@6631.4]
  assign _GEN_939 = {{1'd0}, _T_7190}; // @[Bitwise.scala 48:55:@6632.4]
  assign _T_7242 = _GEN_939 + _T_7241; // @[Bitwise.scala 48:55:@6632.4]
  assign _T_7243 = _T_7193 + _T_7194; // @[Bitwise.scala 48:55:@6633.4]
  assign _T_7244 = _T_7195 + _T_7196; // @[Bitwise.scala 48:55:@6634.4]
  assign _T_7245 = _T_7243 + _T_7244; // @[Bitwise.scala 48:55:@6635.4]
  assign _T_7246 = _T_7242 + _T_7245; // @[Bitwise.scala 48:55:@6636.4]
  assign _T_7247 = _T_7240 + _T_7246; // @[Bitwise.scala 48:55:@6637.4]
  assign _T_7248 = _T_7198 + _T_7199; // @[Bitwise.scala 48:55:@6638.4]
  assign _GEN_940 = {{1'd0}, _T_7197}; // @[Bitwise.scala 48:55:@6639.4]
  assign _T_7249 = _GEN_940 + _T_7248; // @[Bitwise.scala 48:55:@6639.4]
  assign _T_7250 = _T_7200 + _T_7201; // @[Bitwise.scala 48:55:@6640.4]
  assign _T_7251 = _T_7202 + _T_7203; // @[Bitwise.scala 48:55:@6641.4]
  assign _T_7252 = _T_7250 + _T_7251; // @[Bitwise.scala 48:55:@6642.4]
  assign _T_7253 = _T_7249 + _T_7252; // @[Bitwise.scala 48:55:@6643.4]
  assign _T_7254 = _T_7205 + _T_7206; // @[Bitwise.scala 48:55:@6644.4]
  assign _GEN_941 = {{1'd0}, _T_7204}; // @[Bitwise.scala 48:55:@6645.4]
  assign _T_7255 = _GEN_941 + _T_7254; // @[Bitwise.scala 48:55:@6645.4]
  assign _T_7256 = _T_7207 + _T_7208; // @[Bitwise.scala 48:55:@6646.4]
  assign _T_7257 = _T_7209 + _T_7210; // @[Bitwise.scala 48:55:@6647.4]
  assign _T_7258 = _T_7256 + _T_7257; // @[Bitwise.scala 48:55:@6648.4]
  assign _T_7259 = _T_7255 + _T_7258; // @[Bitwise.scala 48:55:@6649.4]
  assign _T_7260 = _T_7253 + _T_7259; // @[Bitwise.scala 48:55:@6650.4]
  assign _T_7261 = _T_7247 + _T_7260; // @[Bitwise.scala 48:55:@6651.4]
  assign _T_7262 = _T_7235 + _T_7261; // @[Bitwise.scala 48:55:@6652.4]
  assign _T_7326 = _T_1124[53:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6717.4]
  assign _T_7327 = _T_7326[0]; // @[Bitwise.scala 50:65:@6718.4]
  assign _T_7328 = _T_7326[1]; // @[Bitwise.scala 50:65:@6719.4]
  assign _T_7329 = _T_7326[2]; // @[Bitwise.scala 50:65:@6720.4]
  assign _T_7330 = _T_7326[3]; // @[Bitwise.scala 50:65:@6721.4]
  assign _T_7331 = _T_7326[4]; // @[Bitwise.scala 50:65:@6722.4]
  assign _T_7332 = _T_7326[5]; // @[Bitwise.scala 50:65:@6723.4]
  assign _T_7333 = _T_7326[6]; // @[Bitwise.scala 50:65:@6724.4]
  assign _T_7334 = _T_7326[7]; // @[Bitwise.scala 50:65:@6725.4]
  assign _T_7335 = _T_7326[8]; // @[Bitwise.scala 50:65:@6726.4]
  assign _T_7336 = _T_7326[9]; // @[Bitwise.scala 50:65:@6727.4]
  assign _T_7337 = _T_7326[10]; // @[Bitwise.scala 50:65:@6728.4]
  assign _T_7338 = _T_7326[11]; // @[Bitwise.scala 50:65:@6729.4]
  assign _T_7339 = _T_7326[12]; // @[Bitwise.scala 50:65:@6730.4]
  assign _T_7340 = _T_7326[13]; // @[Bitwise.scala 50:65:@6731.4]
  assign _T_7341 = _T_7326[14]; // @[Bitwise.scala 50:65:@6732.4]
  assign _T_7342 = _T_7326[15]; // @[Bitwise.scala 50:65:@6733.4]
  assign _T_7343 = _T_7326[16]; // @[Bitwise.scala 50:65:@6734.4]
  assign _T_7344 = _T_7326[17]; // @[Bitwise.scala 50:65:@6735.4]
  assign _T_7345 = _T_7326[18]; // @[Bitwise.scala 50:65:@6736.4]
  assign _T_7346 = _T_7326[19]; // @[Bitwise.scala 50:65:@6737.4]
  assign _T_7347 = _T_7326[20]; // @[Bitwise.scala 50:65:@6738.4]
  assign _T_7348 = _T_7326[21]; // @[Bitwise.scala 50:65:@6739.4]
  assign _T_7349 = _T_7326[22]; // @[Bitwise.scala 50:65:@6740.4]
  assign _T_7350 = _T_7326[23]; // @[Bitwise.scala 50:65:@6741.4]
  assign _T_7351 = _T_7326[24]; // @[Bitwise.scala 50:65:@6742.4]
  assign _T_7352 = _T_7326[25]; // @[Bitwise.scala 50:65:@6743.4]
  assign _T_7353 = _T_7326[26]; // @[Bitwise.scala 50:65:@6744.4]
  assign _T_7354 = _T_7326[27]; // @[Bitwise.scala 50:65:@6745.4]
  assign _T_7355 = _T_7326[28]; // @[Bitwise.scala 50:65:@6746.4]
  assign _T_7356 = _T_7326[29]; // @[Bitwise.scala 50:65:@6747.4]
  assign _T_7357 = _T_7326[30]; // @[Bitwise.scala 50:65:@6748.4]
  assign _T_7358 = _T_7326[31]; // @[Bitwise.scala 50:65:@6749.4]
  assign _T_7359 = _T_7326[32]; // @[Bitwise.scala 50:65:@6750.4]
  assign _T_7360 = _T_7326[33]; // @[Bitwise.scala 50:65:@6751.4]
  assign _T_7361 = _T_7326[34]; // @[Bitwise.scala 50:65:@6752.4]
  assign _T_7362 = _T_7326[35]; // @[Bitwise.scala 50:65:@6753.4]
  assign _T_7363 = _T_7326[36]; // @[Bitwise.scala 50:65:@6754.4]
  assign _T_7364 = _T_7326[37]; // @[Bitwise.scala 50:65:@6755.4]
  assign _T_7365 = _T_7326[38]; // @[Bitwise.scala 50:65:@6756.4]
  assign _T_7366 = _T_7326[39]; // @[Bitwise.scala 50:65:@6757.4]
  assign _T_7367 = _T_7326[40]; // @[Bitwise.scala 50:65:@6758.4]
  assign _T_7368 = _T_7326[41]; // @[Bitwise.scala 50:65:@6759.4]
  assign _T_7369 = _T_7326[42]; // @[Bitwise.scala 50:65:@6760.4]
  assign _T_7370 = _T_7326[43]; // @[Bitwise.scala 50:65:@6761.4]
  assign _T_7371 = _T_7326[44]; // @[Bitwise.scala 50:65:@6762.4]
  assign _T_7372 = _T_7326[45]; // @[Bitwise.scala 50:65:@6763.4]
  assign _T_7373 = _T_7326[46]; // @[Bitwise.scala 50:65:@6764.4]
  assign _T_7374 = _T_7326[47]; // @[Bitwise.scala 50:65:@6765.4]
  assign _T_7375 = _T_7326[48]; // @[Bitwise.scala 50:65:@6766.4]
  assign _T_7376 = _T_7326[49]; // @[Bitwise.scala 50:65:@6767.4]
  assign _T_7377 = _T_7326[50]; // @[Bitwise.scala 50:65:@6768.4]
  assign _T_7378 = _T_7326[51]; // @[Bitwise.scala 50:65:@6769.4]
  assign _T_7379 = _T_7326[52]; // @[Bitwise.scala 50:65:@6770.4]
  assign _T_7380 = _T_7326[53]; // @[Bitwise.scala 50:65:@6771.4]
  assign _T_7381 = _T_7328 + _T_7329; // @[Bitwise.scala 48:55:@6772.4]
  assign _GEN_942 = {{1'd0}, _T_7327}; // @[Bitwise.scala 48:55:@6773.4]
  assign _T_7382 = _GEN_942 + _T_7381; // @[Bitwise.scala 48:55:@6773.4]
  assign _T_7383 = _T_7331 + _T_7332; // @[Bitwise.scala 48:55:@6774.4]
  assign _GEN_943 = {{1'd0}, _T_7330}; // @[Bitwise.scala 48:55:@6775.4]
  assign _T_7384 = _GEN_943 + _T_7383; // @[Bitwise.scala 48:55:@6775.4]
  assign _T_7385 = _T_7382 + _T_7384; // @[Bitwise.scala 48:55:@6776.4]
  assign _T_7386 = _T_7334 + _T_7335; // @[Bitwise.scala 48:55:@6777.4]
  assign _GEN_944 = {{1'd0}, _T_7333}; // @[Bitwise.scala 48:55:@6778.4]
  assign _T_7387 = _GEN_944 + _T_7386; // @[Bitwise.scala 48:55:@6778.4]
  assign _T_7388 = _T_7336 + _T_7337; // @[Bitwise.scala 48:55:@6779.4]
  assign _T_7389 = _T_7338 + _T_7339; // @[Bitwise.scala 48:55:@6780.4]
  assign _T_7390 = _T_7388 + _T_7389; // @[Bitwise.scala 48:55:@6781.4]
  assign _T_7391 = _T_7387 + _T_7390; // @[Bitwise.scala 48:55:@6782.4]
  assign _T_7392 = _T_7385 + _T_7391; // @[Bitwise.scala 48:55:@6783.4]
  assign _T_7393 = _T_7341 + _T_7342; // @[Bitwise.scala 48:55:@6784.4]
  assign _GEN_945 = {{1'd0}, _T_7340}; // @[Bitwise.scala 48:55:@6785.4]
  assign _T_7394 = _GEN_945 + _T_7393; // @[Bitwise.scala 48:55:@6785.4]
  assign _T_7395 = _T_7343 + _T_7344; // @[Bitwise.scala 48:55:@6786.4]
  assign _T_7396 = _T_7345 + _T_7346; // @[Bitwise.scala 48:55:@6787.4]
  assign _T_7397 = _T_7395 + _T_7396; // @[Bitwise.scala 48:55:@6788.4]
  assign _T_7398 = _T_7394 + _T_7397; // @[Bitwise.scala 48:55:@6789.4]
  assign _T_7399 = _T_7348 + _T_7349; // @[Bitwise.scala 48:55:@6790.4]
  assign _GEN_946 = {{1'd0}, _T_7347}; // @[Bitwise.scala 48:55:@6791.4]
  assign _T_7400 = _GEN_946 + _T_7399; // @[Bitwise.scala 48:55:@6791.4]
  assign _T_7401 = _T_7350 + _T_7351; // @[Bitwise.scala 48:55:@6792.4]
  assign _T_7402 = _T_7352 + _T_7353; // @[Bitwise.scala 48:55:@6793.4]
  assign _T_7403 = _T_7401 + _T_7402; // @[Bitwise.scala 48:55:@6794.4]
  assign _T_7404 = _T_7400 + _T_7403; // @[Bitwise.scala 48:55:@6795.4]
  assign _T_7405 = _T_7398 + _T_7404; // @[Bitwise.scala 48:55:@6796.4]
  assign _T_7406 = _T_7392 + _T_7405; // @[Bitwise.scala 48:55:@6797.4]
  assign _T_7407 = _T_7355 + _T_7356; // @[Bitwise.scala 48:55:@6798.4]
  assign _GEN_947 = {{1'd0}, _T_7354}; // @[Bitwise.scala 48:55:@6799.4]
  assign _T_7408 = _GEN_947 + _T_7407; // @[Bitwise.scala 48:55:@6799.4]
  assign _T_7409 = _T_7358 + _T_7359; // @[Bitwise.scala 48:55:@6800.4]
  assign _GEN_948 = {{1'd0}, _T_7357}; // @[Bitwise.scala 48:55:@6801.4]
  assign _T_7410 = _GEN_948 + _T_7409; // @[Bitwise.scala 48:55:@6801.4]
  assign _T_7411 = _T_7408 + _T_7410; // @[Bitwise.scala 48:55:@6802.4]
  assign _T_7412 = _T_7361 + _T_7362; // @[Bitwise.scala 48:55:@6803.4]
  assign _GEN_949 = {{1'd0}, _T_7360}; // @[Bitwise.scala 48:55:@6804.4]
  assign _T_7413 = _GEN_949 + _T_7412; // @[Bitwise.scala 48:55:@6804.4]
  assign _T_7414 = _T_7363 + _T_7364; // @[Bitwise.scala 48:55:@6805.4]
  assign _T_7415 = _T_7365 + _T_7366; // @[Bitwise.scala 48:55:@6806.4]
  assign _T_7416 = _T_7414 + _T_7415; // @[Bitwise.scala 48:55:@6807.4]
  assign _T_7417 = _T_7413 + _T_7416; // @[Bitwise.scala 48:55:@6808.4]
  assign _T_7418 = _T_7411 + _T_7417; // @[Bitwise.scala 48:55:@6809.4]
  assign _T_7419 = _T_7368 + _T_7369; // @[Bitwise.scala 48:55:@6810.4]
  assign _GEN_950 = {{1'd0}, _T_7367}; // @[Bitwise.scala 48:55:@6811.4]
  assign _T_7420 = _GEN_950 + _T_7419; // @[Bitwise.scala 48:55:@6811.4]
  assign _T_7421 = _T_7370 + _T_7371; // @[Bitwise.scala 48:55:@6812.4]
  assign _T_7422 = _T_7372 + _T_7373; // @[Bitwise.scala 48:55:@6813.4]
  assign _T_7423 = _T_7421 + _T_7422; // @[Bitwise.scala 48:55:@6814.4]
  assign _T_7424 = _T_7420 + _T_7423; // @[Bitwise.scala 48:55:@6815.4]
  assign _T_7425 = _T_7375 + _T_7376; // @[Bitwise.scala 48:55:@6816.4]
  assign _GEN_951 = {{1'd0}, _T_7374}; // @[Bitwise.scala 48:55:@6817.4]
  assign _T_7426 = _GEN_951 + _T_7425; // @[Bitwise.scala 48:55:@6817.4]
  assign _T_7427 = _T_7377 + _T_7378; // @[Bitwise.scala 48:55:@6818.4]
  assign _T_7428 = _T_7379 + _T_7380; // @[Bitwise.scala 48:55:@6819.4]
  assign _T_7429 = _T_7427 + _T_7428; // @[Bitwise.scala 48:55:@6820.4]
  assign _T_7430 = _T_7426 + _T_7429; // @[Bitwise.scala 48:55:@6821.4]
  assign _T_7431 = _T_7424 + _T_7430; // @[Bitwise.scala 48:55:@6822.4]
  assign _T_7432 = _T_7418 + _T_7431; // @[Bitwise.scala 48:55:@6823.4]
  assign _T_7433 = _T_7406 + _T_7432; // @[Bitwise.scala 48:55:@6824.4]
  assign _T_7497 = _T_1124[54:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@6889.4]
  assign _T_7498 = _T_7497[0]; // @[Bitwise.scala 50:65:@6890.4]
  assign _T_7499 = _T_7497[1]; // @[Bitwise.scala 50:65:@6891.4]
  assign _T_7500 = _T_7497[2]; // @[Bitwise.scala 50:65:@6892.4]
  assign _T_7501 = _T_7497[3]; // @[Bitwise.scala 50:65:@6893.4]
  assign _T_7502 = _T_7497[4]; // @[Bitwise.scala 50:65:@6894.4]
  assign _T_7503 = _T_7497[5]; // @[Bitwise.scala 50:65:@6895.4]
  assign _T_7504 = _T_7497[6]; // @[Bitwise.scala 50:65:@6896.4]
  assign _T_7505 = _T_7497[7]; // @[Bitwise.scala 50:65:@6897.4]
  assign _T_7506 = _T_7497[8]; // @[Bitwise.scala 50:65:@6898.4]
  assign _T_7507 = _T_7497[9]; // @[Bitwise.scala 50:65:@6899.4]
  assign _T_7508 = _T_7497[10]; // @[Bitwise.scala 50:65:@6900.4]
  assign _T_7509 = _T_7497[11]; // @[Bitwise.scala 50:65:@6901.4]
  assign _T_7510 = _T_7497[12]; // @[Bitwise.scala 50:65:@6902.4]
  assign _T_7511 = _T_7497[13]; // @[Bitwise.scala 50:65:@6903.4]
  assign _T_7512 = _T_7497[14]; // @[Bitwise.scala 50:65:@6904.4]
  assign _T_7513 = _T_7497[15]; // @[Bitwise.scala 50:65:@6905.4]
  assign _T_7514 = _T_7497[16]; // @[Bitwise.scala 50:65:@6906.4]
  assign _T_7515 = _T_7497[17]; // @[Bitwise.scala 50:65:@6907.4]
  assign _T_7516 = _T_7497[18]; // @[Bitwise.scala 50:65:@6908.4]
  assign _T_7517 = _T_7497[19]; // @[Bitwise.scala 50:65:@6909.4]
  assign _T_7518 = _T_7497[20]; // @[Bitwise.scala 50:65:@6910.4]
  assign _T_7519 = _T_7497[21]; // @[Bitwise.scala 50:65:@6911.4]
  assign _T_7520 = _T_7497[22]; // @[Bitwise.scala 50:65:@6912.4]
  assign _T_7521 = _T_7497[23]; // @[Bitwise.scala 50:65:@6913.4]
  assign _T_7522 = _T_7497[24]; // @[Bitwise.scala 50:65:@6914.4]
  assign _T_7523 = _T_7497[25]; // @[Bitwise.scala 50:65:@6915.4]
  assign _T_7524 = _T_7497[26]; // @[Bitwise.scala 50:65:@6916.4]
  assign _T_7525 = _T_7497[27]; // @[Bitwise.scala 50:65:@6917.4]
  assign _T_7526 = _T_7497[28]; // @[Bitwise.scala 50:65:@6918.4]
  assign _T_7527 = _T_7497[29]; // @[Bitwise.scala 50:65:@6919.4]
  assign _T_7528 = _T_7497[30]; // @[Bitwise.scala 50:65:@6920.4]
  assign _T_7529 = _T_7497[31]; // @[Bitwise.scala 50:65:@6921.4]
  assign _T_7530 = _T_7497[32]; // @[Bitwise.scala 50:65:@6922.4]
  assign _T_7531 = _T_7497[33]; // @[Bitwise.scala 50:65:@6923.4]
  assign _T_7532 = _T_7497[34]; // @[Bitwise.scala 50:65:@6924.4]
  assign _T_7533 = _T_7497[35]; // @[Bitwise.scala 50:65:@6925.4]
  assign _T_7534 = _T_7497[36]; // @[Bitwise.scala 50:65:@6926.4]
  assign _T_7535 = _T_7497[37]; // @[Bitwise.scala 50:65:@6927.4]
  assign _T_7536 = _T_7497[38]; // @[Bitwise.scala 50:65:@6928.4]
  assign _T_7537 = _T_7497[39]; // @[Bitwise.scala 50:65:@6929.4]
  assign _T_7538 = _T_7497[40]; // @[Bitwise.scala 50:65:@6930.4]
  assign _T_7539 = _T_7497[41]; // @[Bitwise.scala 50:65:@6931.4]
  assign _T_7540 = _T_7497[42]; // @[Bitwise.scala 50:65:@6932.4]
  assign _T_7541 = _T_7497[43]; // @[Bitwise.scala 50:65:@6933.4]
  assign _T_7542 = _T_7497[44]; // @[Bitwise.scala 50:65:@6934.4]
  assign _T_7543 = _T_7497[45]; // @[Bitwise.scala 50:65:@6935.4]
  assign _T_7544 = _T_7497[46]; // @[Bitwise.scala 50:65:@6936.4]
  assign _T_7545 = _T_7497[47]; // @[Bitwise.scala 50:65:@6937.4]
  assign _T_7546 = _T_7497[48]; // @[Bitwise.scala 50:65:@6938.4]
  assign _T_7547 = _T_7497[49]; // @[Bitwise.scala 50:65:@6939.4]
  assign _T_7548 = _T_7497[50]; // @[Bitwise.scala 50:65:@6940.4]
  assign _T_7549 = _T_7497[51]; // @[Bitwise.scala 50:65:@6941.4]
  assign _T_7550 = _T_7497[52]; // @[Bitwise.scala 50:65:@6942.4]
  assign _T_7551 = _T_7497[53]; // @[Bitwise.scala 50:65:@6943.4]
  assign _T_7552 = _T_7497[54]; // @[Bitwise.scala 50:65:@6944.4]
  assign _T_7553 = _T_7499 + _T_7500; // @[Bitwise.scala 48:55:@6945.4]
  assign _GEN_952 = {{1'd0}, _T_7498}; // @[Bitwise.scala 48:55:@6946.4]
  assign _T_7554 = _GEN_952 + _T_7553; // @[Bitwise.scala 48:55:@6946.4]
  assign _T_7555 = _T_7502 + _T_7503; // @[Bitwise.scala 48:55:@6947.4]
  assign _GEN_953 = {{1'd0}, _T_7501}; // @[Bitwise.scala 48:55:@6948.4]
  assign _T_7556 = _GEN_953 + _T_7555; // @[Bitwise.scala 48:55:@6948.4]
  assign _T_7557 = _T_7554 + _T_7556; // @[Bitwise.scala 48:55:@6949.4]
  assign _T_7558 = _T_7505 + _T_7506; // @[Bitwise.scala 48:55:@6950.4]
  assign _GEN_954 = {{1'd0}, _T_7504}; // @[Bitwise.scala 48:55:@6951.4]
  assign _T_7559 = _GEN_954 + _T_7558; // @[Bitwise.scala 48:55:@6951.4]
  assign _T_7560 = _T_7507 + _T_7508; // @[Bitwise.scala 48:55:@6952.4]
  assign _T_7561 = _T_7509 + _T_7510; // @[Bitwise.scala 48:55:@6953.4]
  assign _T_7562 = _T_7560 + _T_7561; // @[Bitwise.scala 48:55:@6954.4]
  assign _T_7563 = _T_7559 + _T_7562; // @[Bitwise.scala 48:55:@6955.4]
  assign _T_7564 = _T_7557 + _T_7563; // @[Bitwise.scala 48:55:@6956.4]
  assign _T_7565 = _T_7512 + _T_7513; // @[Bitwise.scala 48:55:@6957.4]
  assign _GEN_955 = {{1'd0}, _T_7511}; // @[Bitwise.scala 48:55:@6958.4]
  assign _T_7566 = _GEN_955 + _T_7565; // @[Bitwise.scala 48:55:@6958.4]
  assign _T_7567 = _T_7514 + _T_7515; // @[Bitwise.scala 48:55:@6959.4]
  assign _T_7568 = _T_7516 + _T_7517; // @[Bitwise.scala 48:55:@6960.4]
  assign _T_7569 = _T_7567 + _T_7568; // @[Bitwise.scala 48:55:@6961.4]
  assign _T_7570 = _T_7566 + _T_7569; // @[Bitwise.scala 48:55:@6962.4]
  assign _T_7571 = _T_7519 + _T_7520; // @[Bitwise.scala 48:55:@6963.4]
  assign _GEN_956 = {{1'd0}, _T_7518}; // @[Bitwise.scala 48:55:@6964.4]
  assign _T_7572 = _GEN_956 + _T_7571; // @[Bitwise.scala 48:55:@6964.4]
  assign _T_7573 = _T_7521 + _T_7522; // @[Bitwise.scala 48:55:@6965.4]
  assign _T_7574 = _T_7523 + _T_7524; // @[Bitwise.scala 48:55:@6966.4]
  assign _T_7575 = _T_7573 + _T_7574; // @[Bitwise.scala 48:55:@6967.4]
  assign _T_7576 = _T_7572 + _T_7575; // @[Bitwise.scala 48:55:@6968.4]
  assign _T_7577 = _T_7570 + _T_7576; // @[Bitwise.scala 48:55:@6969.4]
  assign _T_7578 = _T_7564 + _T_7577; // @[Bitwise.scala 48:55:@6970.4]
  assign _T_7579 = _T_7526 + _T_7527; // @[Bitwise.scala 48:55:@6971.4]
  assign _GEN_957 = {{1'd0}, _T_7525}; // @[Bitwise.scala 48:55:@6972.4]
  assign _T_7580 = _GEN_957 + _T_7579; // @[Bitwise.scala 48:55:@6972.4]
  assign _T_7581 = _T_7528 + _T_7529; // @[Bitwise.scala 48:55:@6973.4]
  assign _T_7582 = _T_7530 + _T_7531; // @[Bitwise.scala 48:55:@6974.4]
  assign _T_7583 = _T_7581 + _T_7582; // @[Bitwise.scala 48:55:@6975.4]
  assign _T_7584 = _T_7580 + _T_7583; // @[Bitwise.scala 48:55:@6976.4]
  assign _T_7585 = _T_7533 + _T_7534; // @[Bitwise.scala 48:55:@6977.4]
  assign _GEN_958 = {{1'd0}, _T_7532}; // @[Bitwise.scala 48:55:@6978.4]
  assign _T_7586 = _GEN_958 + _T_7585; // @[Bitwise.scala 48:55:@6978.4]
  assign _T_7587 = _T_7535 + _T_7536; // @[Bitwise.scala 48:55:@6979.4]
  assign _T_7588 = _T_7537 + _T_7538; // @[Bitwise.scala 48:55:@6980.4]
  assign _T_7589 = _T_7587 + _T_7588; // @[Bitwise.scala 48:55:@6981.4]
  assign _T_7590 = _T_7586 + _T_7589; // @[Bitwise.scala 48:55:@6982.4]
  assign _T_7591 = _T_7584 + _T_7590; // @[Bitwise.scala 48:55:@6983.4]
  assign _T_7592 = _T_7540 + _T_7541; // @[Bitwise.scala 48:55:@6984.4]
  assign _GEN_959 = {{1'd0}, _T_7539}; // @[Bitwise.scala 48:55:@6985.4]
  assign _T_7593 = _GEN_959 + _T_7592; // @[Bitwise.scala 48:55:@6985.4]
  assign _T_7594 = _T_7542 + _T_7543; // @[Bitwise.scala 48:55:@6986.4]
  assign _T_7595 = _T_7544 + _T_7545; // @[Bitwise.scala 48:55:@6987.4]
  assign _T_7596 = _T_7594 + _T_7595; // @[Bitwise.scala 48:55:@6988.4]
  assign _T_7597 = _T_7593 + _T_7596; // @[Bitwise.scala 48:55:@6989.4]
  assign _T_7598 = _T_7547 + _T_7548; // @[Bitwise.scala 48:55:@6990.4]
  assign _GEN_960 = {{1'd0}, _T_7546}; // @[Bitwise.scala 48:55:@6991.4]
  assign _T_7599 = _GEN_960 + _T_7598; // @[Bitwise.scala 48:55:@6991.4]
  assign _T_7600 = _T_7549 + _T_7550; // @[Bitwise.scala 48:55:@6992.4]
  assign _T_7601 = _T_7551 + _T_7552; // @[Bitwise.scala 48:55:@6993.4]
  assign _T_7602 = _T_7600 + _T_7601; // @[Bitwise.scala 48:55:@6994.4]
  assign _T_7603 = _T_7599 + _T_7602; // @[Bitwise.scala 48:55:@6995.4]
  assign _T_7604 = _T_7597 + _T_7603; // @[Bitwise.scala 48:55:@6996.4]
  assign _T_7605 = _T_7591 + _T_7604; // @[Bitwise.scala 48:55:@6997.4]
  assign _T_7606 = _T_7578 + _T_7605; // @[Bitwise.scala 48:55:@6998.4]
  assign _T_7670 = _T_1124[55:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7063.4]
  assign _T_7671 = _T_7670[0]; // @[Bitwise.scala 50:65:@7064.4]
  assign _T_7672 = _T_7670[1]; // @[Bitwise.scala 50:65:@7065.4]
  assign _T_7673 = _T_7670[2]; // @[Bitwise.scala 50:65:@7066.4]
  assign _T_7674 = _T_7670[3]; // @[Bitwise.scala 50:65:@7067.4]
  assign _T_7675 = _T_7670[4]; // @[Bitwise.scala 50:65:@7068.4]
  assign _T_7676 = _T_7670[5]; // @[Bitwise.scala 50:65:@7069.4]
  assign _T_7677 = _T_7670[6]; // @[Bitwise.scala 50:65:@7070.4]
  assign _T_7678 = _T_7670[7]; // @[Bitwise.scala 50:65:@7071.4]
  assign _T_7679 = _T_7670[8]; // @[Bitwise.scala 50:65:@7072.4]
  assign _T_7680 = _T_7670[9]; // @[Bitwise.scala 50:65:@7073.4]
  assign _T_7681 = _T_7670[10]; // @[Bitwise.scala 50:65:@7074.4]
  assign _T_7682 = _T_7670[11]; // @[Bitwise.scala 50:65:@7075.4]
  assign _T_7683 = _T_7670[12]; // @[Bitwise.scala 50:65:@7076.4]
  assign _T_7684 = _T_7670[13]; // @[Bitwise.scala 50:65:@7077.4]
  assign _T_7685 = _T_7670[14]; // @[Bitwise.scala 50:65:@7078.4]
  assign _T_7686 = _T_7670[15]; // @[Bitwise.scala 50:65:@7079.4]
  assign _T_7687 = _T_7670[16]; // @[Bitwise.scala 50:65:@7080.4]
  assign _T_7688 = _T_7670[17]; // @[Bitwise.scala 50:65:@7081.4]
  assign _T_7689 = _T_7670[18]; // @[Bitwise.scala 50:65:@7082.4]
  assign _T_7690 = _T_7670[19]; // @[Bitwise.scala 50:65:@7083.4]
  assign _T_7691 = _T_7670[20]; // @[Bitwise.scala 50:65:@7084.4]
  assign _T_7692 = _T_7670[21]; // @[Bitwise.scala 50:65:@7085.4]
  assign _T_7693 = _T_7670[22]; // @[Bitwise.scala 50:65:@7086.4]
  assign _T_7694 = _T_7670[23]; // @[Bitwise.scala 50:65:@7087.4]
  assign _T_7695 = _T_7670[24]; // @[Bitwise.scala 50:65:@7088.4]
  assign _T_7696 = _T_7670[25]; // @[Bitwise.scala 50:65:@7089.4]
  assign _T_7697 = _T_7670[26]; // @[Bitwise.scala 50:65:@7090.4]
  assign _T_7698 = _T_7670[27]; // @[Bitwise.scala 50:65:@7091.4]
  assign _T_7699 = _T_7670[28]; // @[Bitwise.scala 50:65:@7092.4]
  assign _T_7700 = _T_7670[29]; // @[Bitwise.scala 50:65:@7093.4]
  assign _T_7701 = _T_7670[30]; // @[Bitwise.scala 50:65:@7094.4]
  assign _T_7702 = _T_7670[31]; // @[Bitwise.scala 50:65:@7095.4]
  assign _T_7703 = _T_7670[32]; // @[Bitwise.scala 50:65:@7096.4]
  assign _T_7704 = _T_7670[33]; // @[Bitwise.scala 50:65:@7097.4]
  assign _T_7705 = _T_7670[34]; // @[Bitwise.scala 50:65:@7098.4]
  assign _T_7706 = _T_7670[35]; // @[Bitwise.scala 50:65:@7099.4]
  assign _T_7707 = _T_7670[36]; // @[Bitwise.scala 50:65:@7100.4]
  assign _T_7708 = _T_7670[37]; // @[Bitwise.scala 50:65:@7101.4]
  assign _T_7709 = _T_7670[38]; // @[Bitwise.scala 50:65:@7102.4]
  assign _T_7710 = _T_7670[39]; // @[Bitwise.scala 50:65:@7103.4]
  assign _T_7711 = _T_7670[40]; // @[Bitwise.scala 50:65:@7104.4]
  assign _T_7712 = _T_7670[41]; // @[Bitwise.scala 50:65:@7105.4]
  assign _T_7713 = _T_7670[42]; // @[Bitwise.scala 50:65:@7106.4]
  assign _T_7714 = _T_7670[43]; // @[Bitwise.scala 50:65:@7107.4]
  assign _T_7715 = _T_7670[44]; // @[Bitwise.scala 50:65:@7108.4]
  assign _T_7716 = _T_7670[45]; // @[Bitwise.scala 50:65:@7109.4]
  assign _T_7717 = _T_7670[46]; // @[Bitwise.scala 50:65:@7110.4]
  assign _T_7718 = _T_7670[47]; // @[Bitwise.scala 50:65:@7111.4]
  assign _T_7719 = _T_7670[48]; // @[Bitwise.scala 50:65:@7112.4]
  assign _T_7720 = _T_7670[49]; // @[Bitwise.scala 50:65:@7113.4]
  assign _T_7721 = _T_7670[50]; // @[Bitwise.scala 50:65:@7114.4]
  assign _T_7722 = _T_7670[51]; // @[Bitwise.scala 50:65:@7115.4]
  assign _T_7723 = _T_7670[52]; // @[Bitwise.scala 50:65:@7116.4]
  assign _T_7724 = _T_7670[53]; // @[Bitwise.scala 50:65:@7117.4]
  assign _T_7725 = _T_7670[54]; // @[Bitwise.scala 50:65:@7118.4]
  assign _T_7726 = _T_7670[55]; // @[Bitwise.scala 50:65:@7119.4]
  assign _T_7727 = _T_7672 + _T_7673; // @[Bitwise.scala 48:55:@7120.4]
  assign _GEN_961 = {{1'd0}, _T_7671}; // @[Bitwise.scala 48:55:@7121.4]
  assign _T_7728 = _GEN_961 + _T_7727; // @[Bitwise.scala 48:55:@7121.4]
  assign _T_7729 = _T_7674 + _T_7675; // @[Bitwise.scala 48:55:@7122.4]
  assign _T_7730 = _T_7676 + _T_7677; // @[Bitwise.scala 48:55:@7123.4]
  assign _T_7731 = _T_7729 + _T_7730; // @[Bitwise.scala 48:55:@7124.4]
  assign _T_7732 = _T_7728 + _T_7731; // @[Bitwise.scala 48:55:@7125.4]
  assign _T_7733 = _T_7679 + _T_7680; // @[Bitwise.scala 48:55:@7126.4]
  assign _GEN_962 = {{1'd0}, _T_7678}; // @[Bitwise.scala 48:55:@7127.4]
  assign _T_7734 = _GEN_962 + _T_7733; // @[Bitwise.scala 48:55:@7127.4]
  assign _T_7735 = _T_7681 + _T_7682; // @[Bitwise.scala 48:55:@7128.4]
  assign _T_7736 = _T_7683 + _T_7684; // @[Bitwise.scala 48:55:@7129.4]
  assign _T_7737 = _T_7735 + _T_7736; // @[Bitwise.scala 48:55:@7130.4]
  assign _T_7738 = _T_7734 + _T_7737; // @[Bitwise.scala 48:55:@7131.4]
  assign _T_7739 = _T_7732 + _T_7738; // @[Bitwise.scala 48:55:@7132.4]
  assign _T_7740 = _T_7686 + _T_7687; // @[Bitwise.scala 48:55:@7133.4]
  assign _GEN_963 = {{1'd0}, _T_7685}; // @[Bitwise.scala 48:55:@7134.4]
  assign _T_7741 = _GEN_963 + _T_7740; // @[Bitwise.scala 48:55:@7134.4]
  assign _T_7742 = _T_7688 + _T_7689; // @[Bitwise.scala 48:55:@7135.4]
  assign _T_7743 = _T_7690 + _T_7691; // @[Bitwise.scala 48:55:@7136.4]
  assign _T_7744 = _T_7742 + _T_7743; // @[Bitwise.scala 48:55:@7137.4]
  assign _T_7745 = _T_7741 + _T_7744; // @[Bitwise.scala 48:55:@7138.4]
  assign _T_7746 = _T_7693 + _T_7694; // @[Bitwise.scala 48:55:@7139.4]
  assign _GEN_964 = {{1'd0}, _T_7692}; // @[Bitwise.scala 48:55:@7140.4]
  assign _T_7747 = _GEN_964 + _T_7746; // @[Bitwise.scala 48:55:@7140.4]
  assign _T_7748 = _T_7695 + _T_7696; // @[Bitwise.scala 48:55:@7141.4]
  assign _T_7749 = _T_7697 + _T_7698; // @[Bitwise.scala 48:55:@7142.4]
  assign _T_7750 = _T_7748 + _T_7749; // @[Bitwise.scala 48:55:@7143.4]
  assign _T_7751 = _T_7747 + _T_7750; // @[Bitwise.scala 48:55:@7144.4]
  assign _T_7752 = _T_7745 + _T_7751; // @[Bitwise.scala 48:55:@7145.4]
  assign _T_7753 = _T_7739 + _T_7752; // @[Bitwise.scala 48:55:@7146.4]
  assign _T_7754 = _T_7700 + _T_7701; // @[Bitwise.scala 48:55:@7147.4]
  assign _GEN_965 = {{1'd0}, _T_7699}; // @[Bitwise.scala 48:55:@7148.4]
  assign _T_7755 = _GEN_965 + _T_7754; // @[Bitwise.scala 48:55:@7148.4]
  assign _T_7756 = _T_7702 + _T_7703; // @[Bitwise.scala 48:55:@7149.4]
  assign _T_7757 = _T_7704 + _T_7705; // @[Bitwise.scala 48:55:@7150.4]
  assign _T_7758 = _T_7756 + _T_7757; // @[Bitwise.scala 48:55:@7151.4]
  assign _T_7759 = _T_7755 + _T_7758; // @[Bitwise.scala 48:55:@7152.4]
  assign _T_7760 = _T_7707 + _T_7708; // @[Bitwise.scala 48:55:@7153.4]
  assign _GEN_966 = {{1'd0}, _T_7706}; // @[Bitwise.scala 48:55:@7154.4]
  assign _T_7761 = _GEN_966 + _T_7760; // @[Bitwise.scala 48:55:@7154.4]
  assign _T_7762 = _T_7709 + _T_7710; // @[Bitwise.scala 48:55:@7155.4]
  assign _T_7763 = _T_7711 + _T_7712; // @[Bitwise.scala 48:55:@7156.4]
  assign _T_7764 = _T_7762 + _T_7763; // @[Bitwise.scala 48:55:@7157.4]
  assign _T_7765 = _T_7761 + _T_7764; // @[Bitwise.scala 48:55:@7158.4]
  assign _T_7766 = _T_7759 + _T_7765; // @[Bitwise.scala 48:55:@7159.4]
  assign _T_7767 = _T_7714 + _T_7715; // @[Bitwise.scala 48:55:@7160.4]
  assign _GEN_967 = {{1'd0}, _T_7713}; // @[Bitwise.scala 48:55:@7161.4]
  assign _T_7768 = _GEN_967 + _T_7767; // @[Bitwise.scala 48:55:@7161.4]
  assign _T_7769 = _T_7716 + _T_7717; // @[Bitwise.scala 48:55:@7162.4]
  assign _T_7770 = _T_7718 + _T_7719; // @[Bitwise.scala 48:55:@7163.4]
  assign _T_7771 = _T_7769 + _T_7770; // @[Bitwise.scala 48:55:@7164.4]
  assign _T_7772 = _T_7768 + _T_7771; // @[Bitwise.scala 48:55:@7165.4]
  assign _T_7773 = _T_7721 + _T_7722; // @[Bitwise.scala 48:55:@7166.4]
  assign _GEN_968 = {{1'd0}, _T_7720}; // @[Bitwise.scala 48:55:@7167.4]
  assign _T_7774 = _GEN_968 + _T_7773; // @[Bitwise.scala 48:55:@7167.4]
  assign _T_7775 = _T_7723 + _T_7724; // @[Bitwise.scala 48:55:@7168.4]
  assign _T_7776 = _T_7725 + _T_7726; // @[Bitwise.scala 48:55:@7169.4]
  assign _T_7777 = _T_7775 + _T_7776; // @[Bitwise.scala 48:55:@7170.4]
  assign _T_7778 = _T_7774 + _T_7777; // @[Bitwise.scala 48:55:@7171.4]
  assign _T_7779 = _T_7772 + _T_7778; // @[Bitwise.scala 48:55:@7172.4]
  assign _T_7780 = _T_7766 + _T_7779; // @[Bitwise.scala 48:55:@7173.4]
  assign _T_7781 = _T_7753 + _T_7780; // @[Bitwise.scala 48:55:@7174.4]
  assign _T_7845 = _T_1124[56:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7239.4]
  assign _T_7846 = _T_7845[0]; // @[Bitwise.scala 50:65:@7240.4]
  assign _T_7847 = _T_7845[1]; // @[Bitwise.scala 50:65:@7241.4]
  assign _T_7848 = _T_7845[2]; // @[Bitwise.scala 50:65:@7242.4]
  assign _T_7849 = _T_7845[3]; // @[Bitwise.scala 50:65:@7243.4]
  assign _T_7850 = _T_7845[4]; // @[Bitwise.scala 50:65:@7244.4]
  assign _T_7851 = _T_7845[5]; // @[Bitwise.scala 50:65:@7245.4]
  assign _T_7852 = _T_7845[6]; // @[Bitwise.scala 50:65:@7246.4]
  assign _T_7853 = _T_7845[7]; // @[Bitwise.scala 50:65:@7247.4]
  assign _T_7854 = _T_7845[8]; // @[Bitwise.scala 50:65:@7248.4]
  assign _T_7855 = _T_7845[9]; // @[Bitwise.scala 50:65:@7249.4]
  assign _T_7856 = _T_7845[10]; // @[Bitwise.scala 50:65:@7250.4]
  assign _T_7857 = _T_7845[11]; // @[Bitwise.scala 50:65:@7251.4]
  assign _T_7858 = _T_7845[12]; // @[Bitwise.scala 50:65:@7252.4]
  assign _T_7859 = _T_7845[13]; // @[Bitwise.scala 50:65:@7253.4]
  assign _T_7860 = _T_7845[14]; // @[Bitwise.scala 50:65:@7254.4]
  assign _T_7861 = _T_7845[15]; // @[Bitwise.scala 50:65:@7255.4]
  assign _T_7862 = _T_7845[16]; // @[Bitwise.scala 50:65:@7256.4]
  assign _T_7863 = _T_7845[17]; // @[Bitwise.scala 50:65:@7257.4]
  assign _T_7864 = _T_7845[18]; // @[Bitwise.scala 50:65:@7258.4]
  assign _T_7865 = _T_7845[19]; // @[Bitwise.scala 50:65:@7259.4]
  assign _T_7866 = _T_7845[20]; // @[Bitwise.scala 50:65:@7260.4]
  assign _T_7867 = _T_7845[21]; // @[Bitwise.scala 50:65:@7261.4]
  assign _T_7868 = _T_7845[22]; // @[Bitwise.scala 50:65:@7262.4]
  assign _T_7869 = _T_7845[23]; // @[Bitwise.scala 50:65:@7263.4]
  assign _T_7870 = _T_7845[24]; // @[Bitwise.scala 50:65:@7264.4]
  assign _T_7871 = _T_7845[25]; // @[Bitwise.scala 50:65:@7265.4]
  assign _T_7872 = _T_7845[26]; // @[Bitwise.scala 50:65:@7266.4]
  assign _T_7873 = _T_7845[27]; // @[Bitwise.scala 50:65:@7267.4]
  assign _T_7874 = _T_7845[28]; // @[Bitwise.scala 50:65:@7268.4]
  assign _T_7875 = _T_7845[29]; // @[Bitwise.scala 50:65:@7269.4]
  assign _T_7876 = _T_7845[30]; // @[Bitwise.scala 50:65:@7270.4]
  assign _T_7877 = _T_7845[31]; // @[Bitwise.scala 50:65:@7271.4]
  assign _T_7878 = _T_7845[32]; // @[Bitwise.scala 50:65:@7272.4]
  assign _T_7879 = _T_7845[33]; // @[Bitwise.scala 50:65:@7273.4]
  assign _T_7880 = _T_7845[34]; // @[Bitwise.scala 50:65:@7274.4]
  assign _T_7881 = _T_7845[35]; // @[Bitwise.scala 50:65:@7275.4]
  assign _T_7882 = _T_7845[36]; // @[Bitwise.scala 50:65:@7276.4]
  assign _T_7883 = _T_7845[37]; // @[Bitwise.scala 50:65:@7277.4]
  assign _T_7884 = _T_7845[38]; // @[Bitwise.scala 50:65:@7278.4]
  assign _T_7885 = _T_7845[39]; // @[Bitwise.scala 50:65:@7279.4]
  assign _T_7886 = _T_7845[40]; // @[Bitwise.scala 50:65:@7280.4]
  assign _T_7887 = _T_7845[41]; // @[Bitwise.scala 50:65:@7281.4]
  assign _T_7888 = _T_7845[42]; // @[Bitwise.scala 50:65:@7282.4]
  assign _T_7889 = _T_7845[43]; // @[Bitwise.scala 50:65:@7283.4]
  assign _T_7890 = _T_7845[44]; // @[Bitwise.scala 50:65:@7284.4]
  assign _T_7891 = _T_7845[45]; // @[Bitwise.scala 50:65:@7285.4]
  assign _T_7892 = _T_7845[46]; // @[Bitwise.scala 50:65:@7286.4]
  assign _T_7893 = _T_7845[47]; // @[Bitwise.scala 50:65:@7287.4]
  assign _T_7894 = _T_7845[48]; // @[Bitwise.scala 50:65:@7288.4]
  assign _T_7895 = _T_7845[49]; // @[Bitwise.scala 50:65:@7289.4]
  assign _T_7896 = _T_7845[50]; // @[Bitwise.scala 50:65:@7290.4]
  assign _T_7897 = _T_7845[51]; // @[Bitwise.scala 50:65:@7291.4]
  assign _T_7898 = _T_7845[52]; // @[Bitwise.scala 50:65:@7292.4]
  assign _T_7899 = _T_7845[53]; // @[Bitwise.scala 50:65:@7293.4]
  assign _T_7900 = _T_7845[54]; // @[Bitwise.scala 50:65:@7294.4]
  assign _T_7901 = _T_7845[55]; // @[Bitwise.scala 50:65:@7295.4]
  assign _T_7902 = _T_7845[56]; // @[Bitwise.scala 50:65:@7296.4]
  assign _T_7903 = _T_7847 + _T_7848; // @[Bitwise.scala 48:55:@7297.4]
  assign _GEN_969 = {{1'd0}, _T_7846}; // @[Bitwise.scala 48:55:@7298.4]
  assign _T_7904 = _GEN_969 + _T_7903; // @[Bitwise.scala 48:55:@7298.4]
  assign _T_7905 = _T_7849 + _T_7850; // @[Bitwise.scala 48:55:@7299.4]
  assign _T_7906 = _T_7851 + _T_7852; // @[Bitwise.scala 48:55:@7300.4]
  assign _T_7907 = _T_7905 + _T_7906; // @[Bitwise.scala 48:55:@7301.4]
  assign _T_7908 = _T_7904 + _T_7907; // @[Bitwise.scala 48:55:@7302.4]
  assign _T_7909 = _T_7854 + _T_7855; // @[Bitwise.scala 48:55:@7303.4]
  assign _GEN_970 = {{1'd0}, _T_7853}; // @[Bitwise.scala 48:55:@7304.4]
  assign _T_7910 = _GEN_970 + _T_7909; // @[Bitwise.scala 48:55:@7304.4]
  assign _T_7911 = _T_7856 + _T_7857; // @[Bitwise.scala 48:55:@7305.4]
  assign _T_7912 = _T_7858 + _T_7859; // @[Bitwise.scala 48:55:@7306.4]
  assign _T_7913 = _T_7911 + _T_7912; // @[Bitwise.scala 48:55:@7307.4]
  assign _T_7914 = _T_7910 + _T_7913; // @[Bitwise.scala 48:55:@7308.4]
  assign _T_7915 = _T_7908 + _T_7914; // @[Bitwise.scala 48:55:@7309.4]
  assign _T_7916 = _T_7861 + _T_7862; // @[Bitwise.scala 48:55:@7310.4]
  assign _GEN_971 = {{1'd0}, _T_7860}; // @[Bitwise.scala 48:55:@7311.4]
  assign _T_7917 = _GEN_971 + _T_7916; // @[Bitwise.scala 48:55:@7311.4]
  assign _T_7918 = _T_7863 + _T_7864; // @[Bitwise.scala 48:55:@7312.4]
  assign _T_7919 = _T_7865 + _T_7866; // @[Bitwise.scala 48:55:@7313.4]
  assign _T_7920 = _T_7918 + _T_7919; // @[Bitwise.scala 48:55:@7314.4]
  assign _T_7921 = _T_7917 + _T_7920; // @[Bitwise.scala 48:55:@7315.4]
  assign _T_7922 = _T_7868 + _T_7869; // @[Bitwise.scala 48:55:@7316.4]
  assign _GEN_972 = {{1'd0}, _T_7867}; // @[Bitwise.scala 48:55:@7317.4]
  assign _T_7923 = _GEN_972 + _T_7922; // @[Bitwise.scala 48:55:@7317.4]
  assign _T_7924 = _T_7870 + _T_7871; // @[Bitwise.scala 48:55:@7318.4]
  assign _T_7925 = _T_7872 + _T_7873; // @[Bitwise.scala 48:55:@7319.4]
  assign _T_7926 = _T_7924 + _T_7925; // @[Bitwise.scala 48:55:@7320.4]
  assign _T_7927 = _T_7923 + _T_7926; // @[Bitwise.scala 48:55:@7321.4]
  assign _T_7928 = _T_7921 + _T_7927; // @[Bitwise.scala 48:55:@7322.4]
  assign _T_7929 = _T_7915 + _T_7928; // @[Bitwise.scala 48:55:@7323.4]
  assign _T_7930 = _T_7875 + _T_7876; // @[Bitwise.scala 48:55:@7324.4]
  assign _GEN_973 = {{1'd0}, _T_7874}; // @[Bitwise.scala 48:55:@7325.4]
  assign _T_7931 = _GEN_973 + _T_7930; // @[Bitwise.scala 48:55:@7325.4]
  assign _T_7932 = _T_7877 + _T_7878; // @[Bitwise.scala 48:55:@7326.4]
  assign _T_7933 = _T_7879 + _T_7880; // @[Bitwise.scala 48:55:@7327.4]
  assign _T_7934 = _T_7932 + _T_7933; // @[Bitwise.scala 48:55:@7328.4]
  assign _T_7935 = _T_7931 + _T_7934; // @[Bitwise.scala 48:55:@7329.4]
  assign _T_7936 = _T_7882 + _T_7883; // @[Bitwise.scala 48:55:@7330.4]
  assign _GEN_974 = {{1'd0}, _T_7881}; // @[Bitwise.scala 48:55:@7331.4]
  assign _T_7937 = _GEN_974 + _T_7936; // @[Bitwise.scala 48:55:@7331.4]
  assign _T_7938 = _T_7884 + _T_7885; // @[Bitwise.scala 48:55:@7332.4]
  assign _T_7939 = _T_7886 + _T_7887; // @[Bitwise.scala 48:55:@7333.4]
  assign _T_7940 = _T_7938 + _T_7939; // @[Bitwise.scala 48:55:@7334.4]
  assign _T_7941 = _T_7937 + _T_7940; // @[Bitwise.scala 48:55:@7335.4]
  assign _T_7942 = _T_7935 + _T_7941; // @[Bitwise.scala 48:55:@7336.4]
  assign _T_7943 = _T_7889 + _T_7890; // @[Bitwise.scala 48:55:@7337.4]
  assign _GEN_975 = {{1'd0}, _T_7888}; // @[Bitwise.scala 48:55:@7338.4]
  assign _T_7944 = _GEN_975 + _T_7943; // @[Bitwise.scala 48:55:@7338.4]
  assign _T_7945 = _T_7891 + _T_7892; // @[Bitwise.scala 48:55:@7339.4]
  assign _T_7946 = _T_7893 + _T_7894; // @[Bitwise.scala 48:55:@7340.4]
  assign _T_7947 = _T_7945 + _T_7946; // @[Bitwise.scala 48:55:@7341.4]
  assign _T_7948 = _T_7944 + _T_7947; // @[Bitwise.scala 48:55:@7342.4]
  assign _T_7949 = _T_7895 + _T_7896; // @[Bitwise.scala 48:55:@7343.4]
  assign _T_7950 = _T_7897 + _T_7898; // @[Bitwise.scala 48:55:@7344.4]
  assign _T_7951 = _T_7949 + _T_7950; // @[Bitwise.scala 48:55:@7345.4]
  assign _T_7952 = _T_7899 + _T_7900; // @[Bitwise.scala 48:55:@7346.4]
  assign _T_7953 = _T_7901 + _T_7902; // @[Bitwise.scala 48:55:@7347.4]
  assign _T_7954 = _T_7952 + _T_7953; // @[Bitwise.scala 48:55:@7348.4]
  assign _T_7955 = _T_7951 + _T_7954; // @[Bitwise.scala 48:55:@7349.4]
  assign _T_7956 = _T_7948 + _T_7955; // @[Bitwise.scala 48:55:@7350.4]
  assign _T_7957 = _T_7942 + _T_7956; // @[Bitwise.scala 48:55:@7351.4]
  assign _T_7958 = _T_7929 + _T_7957; // @[Bitwise.scala 48:55:@7352.4]
  assign _T_8022 = _T_1124[57:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7417.4]
  assign _T_8023 = _T_8022[0]; // @[Bitwise.scala 50:65:@7418.4]
  assign _T_8024 = _T_8022[1]; // @[Bitwise.scala 50:65:@7419.4]
  assign _T_8025 = _T_8022[2]; // @[Bitwise.scala 50:65:@7420.4]
  assign _T_8026 = _T_8022[3]; // @[Bitwise.scala 50:65:@7421.4]
  assign _T_8027 = _T_8022[4]; // @[Bitwise.scala 50:65:@7422.4]
  assign _T_8028 = _T_8022[5]; // @[Bitwise.scala 50:65:@7423.4]
  assign _T_8029 = _T_8022[6]; // @[Bitwise.scala 50:65:@7424.4]
  assign _T_8030 = _T_8022[7]; // @[Bitwise.scala 50:65:@7425.4]
  assign _T_8031 = _T_8022[8]; // @[Bitwise.scala 50:65:@7426.4]
  assign _T_8032 = _T_8022[9]; // @[Bitwise.scala 50:65:@7427.4]
  assign _T_8033 = _T_8022[10]; // @[Bitwise.scala 50:65:@7428.4]
  assign _T_8034 = _T_8022[11]; // @[Bitwise.scala 50:65:@7429.4]
  assign _T_8035 = _T_8022[12]; // @[Bitwise.scala 50:65:@7430.4]
  assign _T_8036 = _T_8022[13]; // @[Bitwise.scala 50:65:@7431.4]
  assign _T_8037 = _T_8022[14]; // @[Bitwise.scala 50:65:@7432.4]
  assign _T_8038 = _T_8022[15]; // @[Bitwise.scala 50:65:@7433.4]
  assign _T_8039 = _T_8022[16]; // @[Bitwise.scala 50:65:@7434.4]
  assign _T_8040 = _T_8022[17]; // @[Bitwise.scala 50:65:@7435.4]
  assign _T_8041 = _T_8022[18]; // @[Bitwise.scala 50:65:@7436.4]
  assign _T_8042 = _T_8022[19]; // @[Bitwise.scala 50:65:@7437.4]
  assign _T_8043 = _T_8022[20]; // @[Bitwise.scala 50:65:@7438.4]
  assign _T_8044 = _T_8022[21]; // @[Bitwise.scala 50:65:@7439.4]
  assign _T_8045 = _T_8022[22]; // @[Bitwise.scala 50:65:@7440.4]
  assign _T_8046 = _T_8022[23]; // @[Bitwise.scala 50:65:@7441.4]
  assign _T_8047 = _T_8022[24]; // @[Bitwise.scala 50:65:@7442.4]
  assign _T_8048 = _T_8022[25]; // @[Bitwise.scala 50:65:@7443.4]
  assign _T_8049 = _T_8022[26]; // @[Bitwise.scala 50:65:@7444.4]
  assign _T_8050 = _T_8022[27]; // @[Bitwise.scala 50:65:@7445.4]
  assign _T_8051 = _T_8022[28]; // @[Bitwise.scala 50:65:@7446.4]
  assign _T_8052 = _T_8022[29]; // @[Bitwise.scala 50:65:@7447.4]
  assign _T_8053 = _T_8022[30]; // @[Bitwise.scala 50:65:@7448.4]
  assign _T_8054 = _T_8022[31]; // @[Bitwise.scala 50:65:@7449.4]
  assign _T_8055 = _T_8022[32]; // @[Bitwise.scala 50:65:@7450.4]
  assign _T_8056 = _T_8022[33]; // @[Bitwise.scala 50:65:@7451.4]
  assign _T_8057 = _T_8022[34]; // @[Bitwise.scala 50:65:@7452.4]
  assign _T_8058 = _T_8022[35]; // @[Bitwise.scala 50:65:@7453.4]
  assign _T_8059 = _T_8022[36]; // @[Bitwise.scala 50:65:@7454.4]
  assign _T_8060 = _T_8022[37]; // @[Bitwise.scala 50:65:@7455.4]
  assign _T_8061 = _T_8022[38]; // @[Bitwise.scala 50:65:@7456.4]
  assign _T_8062 = _T_8022[39]; // @[Bitwise.scala 50:65:@7457.4]
  assign _T_8063 = _T_8022[40]; // @[Bitwise.scala 50:65:@7458.4]
  assign _T_8064 = _T_8022[41]; // @[Bitwise.scala 50:65:@7459.4]
  assign _T_8065 = _T_8022[42]; // @[Bitwise.scala 50:65:@7460.4]
  assign _T_8066 = _T_8022[43]; // @[Bitwise.scala 50:65:@7461.4]
  assign _T_8067 = _T_8022[44]; // @[Bitwise.scala 50:65:@7462.4]
  assign _T_8068 = _T_8022[45]; // @[Bitwise.scala 50:65:@7463.4]
  assign _T_8069 = _T_8022[46]; // @[Bitwise.scala 50:65:@7464.4]
  assign _T_8070 = _T_8022[47]; // @[Bitwise.scala 50:65:@7465.4]
  assign _T_8071 = _T_8022[48]; // @[Bitwise.scala 50:65:@7466.4]
  assign _T_8072 = _T_8022[49]; // @[Bitwise.scala 50:65:@7467.4]
  assign _T_8073 = _T_8022[50]; // @[Bitwise.scala 50:65:@7468.4]
  assign _T_8074 = _T_8022[51]; // @[Bitwise.scala 50:65:@7469.4]
  assign _T_8075 = _T_8022[52]; // @[Bitwise.scala 50:65:@7470.4]
  assign _T_8076 = _T_8022[53]; // @[Bitwise.scala 50:65:@7471.4]
  assign _T_8077 = _T_8022[54]; // @[Bitwise.scala 50:65:@7472.4]
  assign _T_8078 = _T_8022[55]; // @[Bitwise.scala 50:65:@7473.4]
  assign _T_8079 = _T_8022[56]; // @[Bitwise.scala 50:65:@7474.4]
  assign _T_8080 = _T_8022[57]; // @[Bitwise.scala 50:65:@7475.4]
  assign _T_8081 = _T_8024 + _T_8025; // @[Bitwise.scala 48:55:@7476.4]
  assign _GEN_976 = {{1'd0}, _T_8023}; // @[Bitwise.scala 48:55:@7477.4]
  assign _T_8082 = _GEN_976 + _T_8081; // @[Bitwise.scala 48:55:@7477.4]
  assign _T_8083 = _T_8026 + _T_8027; // @[Bitwise.scala 48:55:@7478.4]
  assign _T_8084 = _T_8028 + _T_8029; // @[Bitwise.scala 48:55:@7479.4]
  assign _T_8085 = _T_8083 + _T_8084; // @[Bitwise.scala 48:55:@7480.4]
  assign _T_8086 = _T_8082 + _T_8085; // @[Bitwise.scala 48:55:@7481.4]
  assign _T_8087 = _T_8031 + _T_8032; // @[Bitwise.scala 48:55:@7482.4]
  assign _GEN_977 = {{1'd0}, _T_8030}; // @[Bitwise.scala 48:55:@7483.4]
  assign _T_8088 = _GEN_977 + _T_8087; // @[Bitwise.scala 48:55:@7483.4]
  assign _T_8089 = _T_8033 + _T_8034; // @[Bitwise.scala 48:55:@7484.4]
  assign _T_8090 = _T_8035 + _T_8036; // @[Bitwise.scala 48:55:@7485.4]
  assign _T_8091 = _T_8089 + _T_8090; // @[Bitwise.scala 48:55:@7486.4]
  assign _T_8092 = _T_8088 + _T_8091; // @[Bitwise.scala 48:55:@7487.4]
  assign _T_8093 = _T_8086 + _T_8092; // @[Bitwise.scala 48:55:@7488.4]
  assign _T_8094 = _T_8038 + _T_8039; // @[Bitwise.scala 48:55:@7489.4]
  assign _GEN_978 = {{1'd0}, _T_8037}; // @[Bitwise.scala 48:55:@7490.4]
  assign _T_8095 = _GEN_978 + _T_8094; // @[Bitwise.scala 48:55:@7490.4]
  assign _T_8096 = _T_8040 + _T_8041; // @[Bitwise.scala 48:55:@7491.4]
  assign _T_8097 = _T_8042 + _T_8043; // @[Bitwise.scala 48:55:@7492.4]
  assign _T_8098 = _T_8096 + _T_8097; // @[Bitwise.scala 48:55:@7493.4]
  assign _T_8099 = _T_8095 + _T_8098; // @[Bitwise.scala 48:55:@7494.4]
  assign _T_8100 = _T_8044 + _T_8045; // @[Bitwise.scala 48:55:@7495.4]
  assign _T_8101 = _T_8046 + _T_8047; // @[Bitwise.scala 48:55:@7496.4]
  assign _T_8102 = _T_8100 + _T_8101; // @[Bitwise.scala 48:55:@7497.4]
  assign _T_8103 = _T_8048 + _T_8049; // @[Bitwise.scala 48:55:@7498.4]
  assign _T_8104 = _T_8050 + _T_8051; // @[Bitwise.scala 48:55:@7499.4]
  assign _T_8105 = _T_8103 + _T_8104; // @[Bitwise.scala 48:55:@7500.4]
  assign _T_8106 = _T_8102 + _T_8105; // @[Bitwise.scala 48:55:@7501.4]
  assign _T_8107 = _T_8099 + _T_8106; // @[Bitwise.scala 48:55:@7502.4]
  assign _T_8108 = _T_8093 + _T_8107; // @[Bitwise.scala 48:55:@7503.4]
  assign _T_8109 = _T_8053 + _T_8054; // @[Bitwise.scala 48:55:@7504.4]
  assign _GEN_979 = {{1'd0}, _T_8052}; // @[Bitwise.scala 48:55:@7505.4]
  assign _T_8110 = _GEN_979 + _T_8109; // @[Bitwise.scala 48:55:@7505.4]
  assign _T_8111 = _T_8055 + _T_8056; // @[Bitwise.scala 48:55:@7506.4]
  assign _T_8112 = _T_8057 + _T_8058; // @[Bitwise.scala 48:55:@7507.4]
  assign _T_8113 = _T_8111 + _T_8112; // @[Bitwise.scala 48:55:@7508.4]
  assign _T_8114 = _T_8110 + _T_8113; // @[Bitwise.scala 48:55:@7509.4]
  assign _T_8115 = _T_8060 + _T_8061; // @[Bitwise.scala 48:55:@7510.4]
  assign _GEN_980 = {{1'd0}, _T_8059}; // @[Bitwise.scala 48:55:@7511.4]
  assign _T_8116 = _GEN_980 + _T_8115; // @[Bitwise.scala 48:55:@7511.4]
  assign _T_8117 = _T_8062 + _T_8063; // @[Bitwise.scala 48:55:@7512.4]
  assign _T_8118 = _T_8064 + _T_8065; // @[Bitwise.scala 48:55:@7513.4]
  assign _T_8119 = _T_8117 + _T_8118; // @[Bitwise.scala 48:55:@7514.4]
  assign _T_8120 = _T_8116 + _T_8119; // @[Bitwise.scala 48:55:@7515.4]
  assign _T_8121 = _T_8114 + _T_8120; // @[Bitwise.scala 48:55:@7516.4]
  assign _T_8122 = _T_8067 + _T_8068; // @[Bitwise.scala 48:55:@7517.4]
  assign _GEN_981 = {{1'd0}, _T_8066}; // @[Bitwise.scala 48:55:@7518.4]
  assign _T_8123 = _GEN_981 + _T_8122; // @[Bitwise.scala 48:55:@7518.4]
  assign _T_8124 = _T_8069 + _T_8070; // @[Bitwise.scala 48:55:@7519.4]
  assign _T_8125 = _T_8071 + _T_8072; // @[Bitwise.scala 48:55:@7520.4]
  assign _T_8126 = _T_8124 + _T_8125; // @[Bitwise.scala 48:55:@7521.4]
  assign _T_8127 = _T_8123 + _T_8126; // @[Bitwise.scala 48:55:@7522.4]
  assign _T_8128 = _T_8073 + _T_8074; // @[Bitwise.scala 48:55:@7523.4]
  assign _T_8129 = _T_8075 + _T_8076; // @[Bitwise.scala 48:55:@7524.4]
  assign _T_8130 = _T_8128 + _T_8129; // @[Bitwise.scala 48:55:@7525.4]
  assign _T_8131 = _T_8077 + _T_8078; // @[Bitwise.scala 48:55:@7526.4]
  assign _T_8132 = _T_8079 + _T_8080; // @[Bitwise.scala 48:55:@7527.4]
  assign _T_8133 = _T_8131 + _T_8132; // @[Bitwise.scala 48:55:@7528.4]
  assign _T_8134 = _T_8130 + _T_8133; // @[Bitwise.scala 48:55:@7529.4]
  assign _T_8135 = _T_8127 + _T_8134; // @[Bitwise.scala 48:55:@7530.4]
  assign _T_8136 = _T_8121 + _T_8135; // @[Bitwise.scala 48:55:@7531.4]
  assign _T_8137 = _T_8108 + _T_8136; // @[Bitwise.scala 48:55:@7532.4]
  assign _T_8201 = _T_1124[58:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7597.4]
  assign _T_8202 = _T_8201[0]; // @[Bitwise.scala 50:65:@7598.4]
  assign _T_8203 = _T_8201[1]; // @[Bitwise.scala 50:65:@7599.4]
  assign _T_8204 = _T_8201[2]; // @[Bitwise.scala 50:65:@7600.4]
  assign _T_8205 = _T_8201[3]; // @[Bitwise.scala 50:65:@7601.4]
  assign _T_8206 = _T_8201[4]; // @[Bitwise.scala 50:65:@7602.4]
  assign _T_8207 = _T_8201[5]; // @[Bitwise.scala 50:65:@7603.4]
  assign _T_8208 = _T_8201[6]; // @[Bitwise.scala 50:65:@7604.4]
  assign _T_8209 = _T_8201[7]; // @[Bitwise.scala 50:65:@7605.4]
  assign _T_8210 = _T_8201[8]; // @[Bitwise.scala 50:65:@7606.4]
  assign _T_8211 = _T_8201[9]; // @[Bitwise.scala 50:65:@7607.4]
  assign _T_8212 = _T_8201[10]; // @[Bitwise.scala 50:65:@7608.4]
  assign _T_8213 = _T_8201[11]; // @[Bitwise.scala 50:65:@7609.4]
  assign _T_8214 = _T_8201[12]; // @[Bitwise.scala 50:65:@7610.4]
  assign _T_8215 = _T_8201[13]; // @[Bitwise.scala 50:65:@7611.4]
  assign _T_8216 = _T_8201[14]; // @[Bitwise.scala 50:65:@7612.4]
  assign _T_8217 = _T_8201[15]; // @[Bitwise.scala 50:65:@7613.4]
  assign _T_8218 = _T_8201[16]; // @[Bitwise.scala 50:65:@7614.4]
  assign _T_8219 = _T_8201[17]; // @[Bitwise.scala 50:65:@7615.4]
  assign _T_8220 = _T_8201[18]; // @[Bitwise.scala 50:65:@7616.4]
  assign _T_8221 = _T_8201[19]; // @[Bitwise.scala 50:65:@7617.4]
  assign _T_8222 = _T_8201[20]; // @[Bitwise.scala 50:65:@7618.4]
  assign _T_8223 = _T_8201[21]; // @[Bitwise.scala 50:65:@7619.4]
  assign _T_8224 = _T_8201[22]; // @[Bitwise.scala 50:65:@7620.4]
  assign _T_8225 = _T_8201[23]; // @[Bitwise.scala 50:65:@7621.4]
  assign _T_8226 = _T_8201[24]; // @[Bitwise.scala 50:65:@7622.4]
  assign _T_8227 = _T_8201[25]; // @[Bitwise.scala 50:65:@7623.4]
  assign _T_8228 = _T_8201[26]; // @[Bitwise.scala 50:65:@7624.4]
  assign _T_8229 = _T_8201[27]; // @[Bitwise.scala 50:65:@7625.4]
  assign _T_8230 = _T_8201[28]; // @[Bitwise.scala 50:65:@7626.4]
  assign _T_8231 = _T_8201[29]; // @[Bitwise.scala 50:65:@7627.4]
  assign _T_8232 = _T_8201[30]; // @[Bitwise.scala 50:65:@7628.4]
  assign _T_8233 = _T_8201[31]; // @[Bitwise.scala 50:65:@7629.4]
  assign _T_8234 = _T_8201[32]; // @[Bitwise.scala 50:65:@7630.4]
  assign _T_8235 = _T_8201[33]; // @[Bitwise.scala 50:65:@7631.4]
  assign _T_8236 = _T_8201[34]; // @[Bitwise.scala 50:65:@7632.4]
  assign _T_8237 = _T_8201[35]; // @[Bitwise.scala 50:65:@7633.4]
  assign _T_8238 = _T_8201[36]; // @[Bitwise.scala 50:65:@7634.4]
  assign _T_8239 = _T_8201[37]; // @[Bitwise.scala 50:65:@7635.4]
  assign _T_8240 = _T_8201[38]; // @[Bitwise.scala 50:65:@7636.4]
  assign _T_8241 = _T_8201[39]; // @[Bitwise.scala 50:65:@7637.4]
  assign _T_8242 = _T_8201[40]; // @[Bitwise.scala 50:65:@7638.4]
  assign _T_8243 = _T_8201[41]; // @[Bitwise.scala 50:65:@7639.4]
  assign _T_8244 = _T_8201[42]; // @[Bitwise.scala 50:65:@7640.4]
  assign _T_8245 = _T_8201[43]; // @[Bitwise.scala 50:65:@7641.4]
  assign _T_8246 = _T_8201[44]; // @[Bitwise.scala 50:65:@7642.4]
  assign _T_8247 = _T_8201[45]; // @[Bitwise.scala 50:65:@7643.4]
  assign _T_8248 = _T_8201[46]; // @[Bitwise.scala 50:65:@7644.4]
  assign _T_8249 = _T_8201[47]; // @[Bitwise.scala 50:65:@7645.4]
  assign _T_8250 = _T_8201[48]; // @[Bitwise.scala 50:65:@7646.4]
  assign _T_8251 = _T_8201[49]; // @[Bitwise.scala 50:65:@7647.4]
  assign _T_8252 = _T_8201[50]; // @[Bitwise.scala 50:65:@7648.4]
  assign _T_8253 = _T_8201[51]; // @[Bitwise.scala 50:65:@7649.4]
  assign _T_8254 = _T_8201[52]; // @[Bitwise.scala 50:65:@7650.4]
  assign _T_8255 = _T_8201[53]; // @[Bitwise.scala 50:65:@7651.4]
  assign _T_8256 = _T_8201[54]; // @[Bitwise.scala 50:65:@7652.4]
  assign _T_8257 = _T_8201[55]; // @[Bitwise.scala 50:65:@7653.4]
  assign _T_8258 = _T_8201[56]; // @[Bitwise.scala 50:65:@7654.4]
  assign _T_8259 = _T_8201[57]; // @[Bitwise.scala 50:65:@7655.4]
  assign _T_8260 = _T_8201[58]; // @[Bitwise.scala 50:65:@7656.4]
  assign _T_8261 = _T_8203 + _T_8204; // @[Bitwise.scala 48:55:@7657.4]
  assign _GEN_982 = {{1'd0}, _T_8202}; // @[Bitwise.scala 48:55:@7658.4]
  assign _T_8262 = _GEN_982 + _T_8261; // @[Bitwise.scala 48:55:@7658.4]
  assign _T_8263 = _T_8205 + _T_8206; // @[Bitwise.scala 48:55:@7659.4]
  assign _T_8264 = _T_8207 + _T_8208; // @[Bitwise.scala 48:55:@7660.4]
  assign _T_8265 = _T_8263 + _T_8264; // @[Bitwise.scala 48:55:@7661.4]
  assign _T_8266 = _T_8262 + _T_8265; // @[Bitwise.scala 48:55:@7662.4]
  assign _T_8267 = _T_8210 + _T_8211; // @[Bitwise.scala 48:55:@7663.4]
  assign _GEN_983 = {{1'd0}, _T_8209}; // @[Bitwise.scala 48:55:@7664.4]
  assign _T_8268 = _GEN_983 + _T_8267; // @[Bitwise.scala 48:55:@7664.4]
  assign _T_8269 = _T_8212 + _T_8213; // @[Bitwise.scala 48:55:@7665.4]
  assign _T_8270 = _T_8214 + _T_8215; // @[Bitwise.scala 48:55:@7666.4]
  assign _T_8271 = _T_8269 + _T_8270; // @[Bitwise.scala 48:55:@7667.4]
  assign _T_8272 = _T_8268 + _T_8271; // @[Bitwise.scala 48:55:@7668.4]
  assign _T_8273 = _T_8266 + _T_8272; // @[Bitwise.scala 48:55:@7669.4]
  assign _T_8274 = _T_8217 + _T_8218; // @[Bitwise.scala 48:55:@7670.4]
  assign _GEN_984 = {{1'd0}, _T_8216}; // @[Bitwise.scala 48:55:@7671.4]
  assign _T_8275 = _GEN_984 + _T_8274; // @[Bitwise.scala 48:55:@7671.4]
  assign _T_8276 = _T_8219 + _T_8220; // @[Bitwise.scala 48:55:@7672.4]
  assign _T_8277 = _T_8221 + _T_8222; // @[Bitwise.scala 48:55:@7673.4]
  assign _T_8278 = _T_8276 + _T_8277; // @[Bitwise.scala 48:55:@7674.4]
  assign _T_8279 = _T_8275 + _T_8278; // @[Bitwise.scala 48:55:@7675.4]
  assign _T_8280 = _T_8223 + _T_8224; // @[Bitwise.scala 48:55:@7676.4]
  assign _T_8281 = _T_8225 + _T_8226; // @[Bitwise.scala 48:55:@7677.4]
  assign _T_8282 = _T_8280 + _T_8281; // @[Bitwise.scala 48:55:@7678.4]
  assign _T_8283 = _T_8227 + _T_8228; // @[Bitwise.scala 48:55:@7679.4]
  assign _T_8284 = _T_8229 + _T_8230; // @[Bitwise.scala 48:55:@7680.4]
  assign _T_8285 = _T_8283 + _T_8284; // @[Bitwise.scala 48:55:@7681.4]
  assign _T_8286 = _T_8282 + _T_8285; // @[Bitwise.scala 48:55:@7682.4]
  assign _T_8287 = _T_8279 + _T_8286; // @[Bitwise.scala 48:55:@7683.4]
  assign _T_8288 = _T_8273 + _T_8287; // @[Bitwise.scala 48:55:@7684.4]
  assign _T_8289 = _T_8232 + _T_8233; // @[Bitwise.scala 48:55:@7685.4]
  assign _GEN_985 = {{1'd0}, _T_8231}; // @[Bitwise.scala 48:55:@7686.4]
  assign _T_8290 = _GEN_985 + _T_8289; // @[Bitwise.scala 48:55:@7686.4]
  assign _T_8291 = _T_8234 + _T_8235; // @[Bitwise.scala 48:55:@7687.4]
  assign _T_8292 = _T_8236 + _T_8237; // @[Bitwise.scala 48:55:@7688.4]
  assign _T_8293 = _T_8291 + _T_8292; // @[Bitwise.scala 48:55:@7689.4]
  assign _T_8294 = _T_8290 + _T_8293; // @[Bitwise.scala 48:55:@7690.4]
  assign _T_8295 = _T_8238 + _T_8239; // @[Bitwise.scala 48:55:@7691.4]
  assign _T_8296 = _T_8240 + _T_8241; // @[Bitwise.scala 48:55:@7692.4]
  assign _T_8297 = _T_8295 + _T_8296; // @[Bitwise.scala 48:55:@7693.4]
  assign _T_8298 = _T_8242 + _T_8243; // @[Bitwise.scala 48:55:@7694.4]
  assign _T_8299 = _T_8244 + _T_8245; // @[Bitwise.scala 48:55:@7695.4]
  assign _T_8300 = _T_8298 + _T_8299; // @[Bitwise.scala 48:55:@7696.4]
  assign _T_8301 = _T_8297 + _T_8300; // @[Bitwise.scala 48:55:@7697.4]
  assign _T_8302 = _T_8294 + _T_8301; // @[Bitwise.scala 48:55:@7698.4]
  assign _T_8303 = _T_8247 + _T_8248; // @[Bitwise.scala 48:55:@7699.4]
  assign _GEN_986 = {{1'd0}, _T_8246}; // @[Bitwise.scala 48:55:@7700.4]
  assign _T_8304 = _GEN_986 + _T_8303; // @[Bitwise.scala 48:55:@7700.4]
  assign _T_8305 = _T_8249 + _T_8250; // @[Bitwise.scala 48:55:@7701.4]
  assign _T_8306 = _T_8251 + _T_8252; // @[Bitwise.scala 48:55:@7702.4]
  assign _T_8307 = _T_8305 + _T_8306; // @[Bitwise.scala 48:55:@7703.4]
  assign _T_8308 = _T_8304 + _T_8307; // @[Bitwise.scala 48:55:@7704.4]
  assign _T_8309 = _T_8253 + _T_8254; // @[Bitwise.scala 48:55:@7705.4]
  assign _T_8310 = _T_8255 + _T_8256; // @[Bitwise.scala 48:55:@7706.4]
  assign _T_8311 = _T_8309 + _T_8310; // @[Bitwise.scala 48:55:@7707.4]
  assign _T_8312 = _T_8257 + _T_8258; // @[Bitwise.scala 48:55:@7708.4]
  assign _T_8313 = _T_8259 + _T_8260; // @[Bitwise.scala 48:55:@7709.4]
  assign _T_8314 = _T_8312 + _T_8313; // @[Bitwise.scala 48:55:@7710.4]
  assign _T_8315 = _T_8311 + _T_8314; // @[Bitwise.scala 48:55:@7711.4]
  assign _T_8316 = _T_8308 + _T_8315; // @[Bitwise.scala 48:55:@7712.4]
  assign _T_8317 = _T_8302 + _T_8316; // @[Bitwise.scala 48:55:@7713.4]
  assign _T_8318 = _T_8288 + _T_8317; // @[Bitwise.scala 48:55:@7714.4]
  assign _T_8382 = _T_1124[59:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7779.4]
  assign _T_8383 = _T_8382[0]; // @[Bitwise.scala 50:65:@7780.4]
  assign _T_8384 = _T_8382[1]; // @[Bitwise.scala 50:65:@7781.4]
  assign _T_8385 = _T_8382[2]; // @[Bitwise.scala 50:65:@7782.4]
  assign _T_8386 = _T_8382[3]; // @[Bitwise.scala 50:65:@7783.4]
  assign _T_8387 = _T_8382[4]; // @[Bitwise.scala 50:65:@7784.4]
  assign _T_8388 = _T_8382[5]; // @[Bitwise.scala 50:65:@7785.4]
  assign _T_8389 = _T_8382[6]; // @[Bitwise.scala 50:65:@7786.4]
  assign _T_8390 = _T_8382[7]; // @[Bitwise.scala 50:65:@7787.4]
  assign _T_8391 = _T_8382[8]; // @[Bitwise.scala 50:65:@7788.4]
  assign _T_8392 = _T_8382[9]; // @[Bitwise.scala 50:65:@7789.4]
  assign _T_8393 = _T_8382[10]; // @[Bitwise.scala 50:65:@7790.4]
  assign _T_8394 = _T_8382[11]; // @[Bitwise.scala 50:65:@7791.4]
  assign _T_8395 = _T_8382[12]; // @[Bitwise.scala 50:65:@7792.4]
  assign _T_8396 = _T_8382[13]; // @[Bitwise.scala 50:65:@7793.4]
  assign _T_8397 = _T_8382[14]; // @[Bitwise.scala 50:65:@7794.4]
  assign _T_8398 = _T_8382[15]; // @[Bitwise.scala 50:65:@7795.4]
  assign _T_8399 = _T_8382[16]; // @[Bitwise.scala 50:65:@7796.4]
  assign _T_8400 = _T_8382[17]; // @[Bitwise.scala 50:65:@7797.4]
  assign _T_8401 = _T_8382[18]; // @[Bitwise.scala 50:65:@7798.4]
  assign _T_8402 = _T_8382[19]; // @[Bitwise.scala 50:65:@7799.4]
  assign _T_8403 = _T_8382[20]; // @[Bitwise.scala 50:65:@7800.4]
  assign _T_8404 = _T_8382[21]; // @[Bitwise.scala 50:65:@7801.4]
  assign _T_8405 = _T_8382[22]; // @[Bitwise.scala 50:65:@7802.4]
  assign _T_8406 = _T_8382[23]; // @[Bitwise.scala 50:65:@7803.4]
  assign _T_8407 = _T_8382[24]; // @[Bitwise.scala 50:65:@7804.4]
  assign _T_8408 = _T_8382[25]; // @[Bitwise.scala 50:65:@7805.4]
  assign _T_8409 = _T_8382[26]; // @[Bitwise.scala 50:65:@7806.4]
  assign _T_8410 = _T_8382[27]; // @[Bitwise.scala 50:65:@7807.4]
  assign _T_8411 = _T_8382[28]; // @[Bitwise.scala 50:65:@7808.4]
  assign _T_8412 = _T_8382[29]; // @[Bitwise.scala 50:65:@7809.4]
  assign _T_8413 = _T_8382[30]; // @[Bitwise.scala 50:65:@7810.4]
  assign _T_8414 = _T_8382[31]; // @[Bitwise.scala 50:65:@7811.4]
  assign _T_8415 = _T_8382[32]; // @[Bitwise.scala 50:65:@7812.4]
  assign _T_8416 = _T_8382[33]; // @[Bitwise.scala 50:65:@7813.4]
  assign _T_8417 = _T_8382[34]; // @[Bitwise.scala 50:65:@7814.4]
  assign _T_8418 = _T_8382[35]; // @[Bitwise.scala 50:65:@7815.4]
  assign _T_8419 = _T_8382[36]; // @[Bitwise.scala 50:65:@7816.4]
  assign _T_8420 = _T_8382[37]; // @[Bitwise.scala 50:65:@7817.4]
  assign _T_8421 = _T_8382[38]; // @[Bitwise.scala 50:65:@7818.4]
  assign _T_8422 = _T_8382[39]; // @[Bitwise.scala 50:65:@7819.4]
  assign _T_8423 = _T_8382[40]; // @[Bitwise.scala 50:65:@7820.4]
  assign _T_8424 = _T_8382[41]; // @[Bitwise.scala 50:65:@7821.4]
  assign _T_8425 = _T_8382[42]; // @[Bitwise.scala 50:65:@7822.4]
  assign _T_8426 = _T_8382[43]; // @[Bitwise.scala 50:65:@7823.4]
  assign _T_8427 = _T_8382[44]; // @[Bitwise.scala 50:65:@7824.4]
  assign _T_8428 = _T_8382[45]; // @[Bitwise.scala 50:65:@7825.4]
  assign _T_8429 = _T_8382[46]; // @[Bitwise.scala 50:65:@7826.4]
  assign _T_8430 = _T_8382[47]; // @[Bitwise.scala 50:65:@7827.4]
  assign _T_8431 = _T_8382[48]; // @[Bitwise.scala 50:65:@7828.4]
  assign _T_8432 = _T_8382[49]; // @[Bitwise.scala 50:65:@7829.4]
  assign _T_8433 = _T_8382[50]; // @[Bitwise.scala 50:65:@7830.4]
  assign _T_8434 = _T_8382[51]; // @[Bitwise.scala 50:65:@7831.4]
  assign _T_8435 = _T_8382[52]; // @[Bitwise.scala 50:65:@7832.4]
  assign _T_8436 = _T_8382[53]; // @[Bitwise.scala 50:65:@7833.4]
  assign _T_8437 = _T_8382[54]; // @[Bitwise.scala 50:65:@7834.4]
  assign _T_8438 = _T_8382[55]; // @[Bitwise.scala 50:65:@7835.4]
  assign _T_8439 = _T_8382[56]; // @[Bitwise.scala 50:65:@7836.4]
  assign _T_8440 = _T_8382[57]; // @[Bitwise.scala 50:65:@7837.4]
  assign _T_8441 = _T_8382[58]; // @[Bitwise.scala 50:65:@7838.4]
  assign _T_8442 = _T_8382[59]; // @[Bitwise.scala 50:65:@7839.4]
  assign _T_8443 = _T_8384 + _T_8385; // @[Bitwise.scala 48:55:@7840.4]
  assign _GEN_987 = {{1'd0}, _T_8383}; // @[Bitwise.scala 48:55:@7841.4]
  assign _T_8444 = _GEN_987 + _T_8443; // @[Bitwise.scala 48:55:@7841.4]
  assign _T_8445 = _T_8386 + _T_8387; // @[Bitwise.scala 48:55:@7842.4]
  assign _T_8446 = _T_8388 + _T_8389; // @[Bitwise.scala 48:55:@7843.4]
  assign _T_8447 = _T_8445 + _T_8446; // @[Bitwise.scala 48:55:@7844.4]
  assign _T_8448 = _T_8444 + _T_8447; // @[Bitwise.scala 48:55:@7845.4]
  assign _T_8449 = _T_8390 + _T_8391; // @[Bitwise.scala 48:55:@7846.4]
  assign _T_8450 = _T_8392 + _T_8393; // @[Bitwise.scala 48:55:@7847.4]
  assign _T_8451 = _T_8449 + _T_8450; // @[Bitwise.scala 48:55:@7848.4]
  assign _T_8452 = _T_8394 + _T_8395; // @[Bitwise.scala 48:55:@7849.4]
  assign _T_8453 = _T_8396 + _T_8397; // @[Bitwise.scala 48:55:@7850.4]
  assign _T_8454 = _T_8452 + _T_8453; // @[Bitwise.scala 48:55:@7851.4]
  assign _T_8455 = _T_8451 + _T_8454; // @[Bitwise.scala 48:55:@7852.4]
  assign _T_8456 = _T_8448 + _T_8455; // @[Bitwise.scala 48:55:@7853.4]
  assign _T_8457 = _T_8399 + _T_8400; // @[Bitwise.scala 48:55:@7854.4]
  assign _GEN_988 = {{1'd0}, _T_8398}; // @[Bitwise.scala 48:55:@7855.4]
  assign _T_8458 = _GEN_988 + _T_8457; // @[Bitwise.scala 48:55:@7855.4]
  assign _T_8459 = _T_8401 + _T_8402; // @[Bitwise.scala 48:55:@7856.4]
  assign _T_8460 = _T_8403 + _T_8404; // @[Bitwise.scala 48:55:@7857.4]
  assign _T_8461 = _T_8459 + _T_8460; // @[Bitwise.scala 48:55:@7858.4]
  assign _T_8462 = _T_8458 + _T_8461; // @[Bitwise.scala 48:55:@7859.4]
  assign _T_8463 = _T_8405 + _T_8406; // @[Bitwise.scala 48:55:@7860.4]
  assign _T_8464 = _T_8407 + _T_8408; // @[Bitwise.scala 48:55:@7861.4]
  assign _T_8465 = _T_8463 + _T_8464; // @[Bitwise.scala 48:55:@7862.4]
  assign _T_8466 = _T_8409 + _T_8410; // @[Bitwise.scala 48:55:@7863.4]
  assign _T_8467 = _T_8411 + _T_8412; // @[Bitwise.scala 48:55:@7864.4]
  assign _T_8468 = _T_8466 + _T_8467; // @[Bitwise.scala 48:55:@7865.4]
  assign _T_8469 = _T_8465 + _T_8468; // @[Bitwise.scala 48:55:@7866.4]
  assign _T_8470 = _T_8462 + _T_8469; // @[Bitwise.scala 48:55:@7867.4]
  assign _T_8471 = _T_8456 + _T_8470; // @[Bitwise.scala 48:55:@7868.4]
  assign _T_8472 = _T_8414 + _T_8415; // @[Bitwise.scala 48:55:@7869.4]
  assign _GEN_989 = {{1'd0}, _T_8413}; // @[Bitwise.scala 48:55:@7870.4]
  assign _T_8473 = _GEN_989 + _T_8472; // @[Bitwise.scala 48:55:@7870.4]
  assign _T_8474 = _T_8416 + _T_8417; // @[Bitwise.scala 48:55:@7871.4]
  assign _T_8475 = _T_8418 + _T_8419; // @[Bitwise.scala 48:55:@7872.4]
  assign _T_8476 = _T_8474 + _T_8475; // @[Bitwise.scala 48:55:@7873.4]
  assign _T_8477 = _T_8473 + _T_8476; // @[Bitwise.scala 48:55:@7874.4]
  assign _T_8478 = _T_8420 + _T_8421; // @[Bitwise.scala 48:55:@7875.4]
  assign _T_8479 = _T_8422 + _T_8423; // @[Bitwise.scala 48:55:@7876.4]
  assign _T_8480 = _T_8478 + _T_8479; // @[Bitwise.scala 48:55:@7877.4]
  assign _T_8481 = _T_8424 + _T_8425; // @[Bitwise.scala 48:55:@7878.4]
  assign _T_8482 = _T_8426 + _T_8427; // @[Bitwise.scala 48:55:@7879.4]
  assign _T_8483 = _T_8481 + _T_8482; // @[Bitwise.scala 48:55:@7880.4]
  assign _T_8484 = _T_8480 + _T_8483; // @[Bitwise.scala 48:55:@7881.4]
  assign _T_8485 = _T_8477 + _T_8484; // @[Bitwise.scala 48:55:@7882.4]
  assign _T_8486 = _T_8429 + _T_8430; // @[Bitwise.scala 48:55:@7883.4]
  assign _GEN_990 = {{1'd0}, _T_8428}; // @[Bitwise.scala 48:55:@7884.4]
  assign _T_8487 = _GEN_990 + _T_8486; // @[Bitwise.scala 48:55:@7884.4]
  assign _T_8488 = _T_8431 + _T_8432; // @[Bitwise.scala 48:55:@7885.4]
  assign _T_8489 = _T_8433 + _T_8434; // @[Bitwise.scala 48:55:@7886.4]
  assign _T_8490 = _T_8488 + _T_8489; // @[Bitwise.scala 48:55:@7887.4]
  assign _T_8491 = _T_8487 + _T_8490; // @[Bitwise.scala 48:55:@7888.4]
  assign _T_8492 = _T_8435 + _T_8436; // @[Bitwise.scala 48:55:@7889.4]
  assign _T_8493 = _T_8437 + _T_8438; // @[Bitwise.scala 48:55:@7890.4]
  assign _T_8494 = _T_8492 + _T_8493; // @[Bitwise.scala 48:55:@7891.4]
  assign _T_8495 = _T_8439 + _T_8440; // @[Bitwise.scala 48:55:@7892.4]
  assign _T_8496 = _T_8441 + _T_8442; // @[Bitwise.scala 48:55:@7893.4]
  assign _T_8497 = _T_8495 + _T_8496; // @[Bitwise.scala 48:55:@7894.4]
  assign _T_8498 = _T_8494 + _T_8497; // @[Bitwise.scala 48:55:@7895.4]
  assign _T_8499 = _T_8491 + _T_8498; // @[Bitwise.scala 48:55:@7896.4]
  assign _T_8500 = _T_8485 + _T_8499; // @[Bitwise.scala 48:55:@7897.4]
  assign _T_8501 = _T_8471 + _T_8500; // @[Bitwise.scala 48:55:@7898.4]
  assign _T_8565 = _T_1124[60:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@7963.4]
  assign _T_8566 = _T_8565[0]; // @[Bitwise.scala 50:65:@7964.4]
  assign _T_8567 = _T_8565[1]; // @[Bitwise.scala 50:65:@7965.4]
  assign _T_8568 = _T_8565[2]; // @[Bitwise.scala 50:65:@7966.4]
  assign _T_8569 = _T_8565[3]; // @[Bitwise.scala 50:65:@7967.4]
  assign _T_8570 = _T_8565[4]; // @[Bitwise.scala 50:65:@7968.4]
  assign _T_8571 = _T_8565[5]; // @[Bitwise.scala 50:65:@7969.4]
  assign _T_8572 = _T_8565[6]; // @[Bitwise.scala 50:65:@7970.4]
  assign _T_8573 = _T_8565[7]; // @[Bitwise.scala 50:65:@7971.4]
  assign _T_8574 = _T_8565[8]; // @[Bitwise.scala 50:65:@7972.4]
  assign _T_8575 = _T_8565[9]; // @[Bitwise.scala 50:65:@7973.4]
  assign _T_8576 = _T_8565[10]; // @[Bitwise.scala 50:65:@7974.4]
  assign _T_8577 = _T_8565[11]; // @[Bitwise.scala 50:65:@7975.4]
  assign _T_8578 = _T_8565[12]; // @[Bitwise.scala 50:65:@7976.4]
  assign _T_8579 = _T_8565[13]; // @[Bitwise.scala 50:65:@7977.4]
  assign _T_8580 = _T_8565[14]; // @[Bitwise.scala 50:65:@7978.4]
  assign _T_8581 = _T_8565[15]; // @[Bitwise.scala 50:65:@7979.4]
  assign _T_8582 = _T_8565[16]; // @[Bitwise.scala 50:65:@7980.4]
  assign _T_8583 = _T_8565[17]; // @[Bitwise.scala 50:65:@7981.4]
  assign _T_8584 = _T_8565[18]; // @[Bitwise.scala 50:65:@7982.4]
  assign _T_8585 = _T_8565[19]; // @[Bitwise.scala 50:65:@7983.4]
  assign _T_8586 = _T_8565[20]; // @[Bitwise.scala 50:65:@7984.4]
  assign _T_8587 = _T_8565[21]; // @[Bitwise.scala 50:65:@7985.4]
  assign _T_8588 = _T_8565[22]; // @[Bitwise.scala 50:65:@7986.4]
  assign _T_8589 = _T_8565[23]; // @[Bitwise.scala 50:65:@7987.4]
  assign _T_8590 = _T_8565[24]; // @[Bitwise.scala 50:65:@7988.4]
  assign _T_8591 = _T_8565[25]; // @[Bitwise.scala 50:65:@7989.4]
  assign _T_8592 = _T_8565[26]; // @[Bitwise.scala 50:65:@7990.4]
  assign _T_8593 = _T_8565[27]; // @[Bitwise.scala 50:65:@7991.4]
  assign _T_8594 = _T_8565[28]; // @[Bitwise.scala 50:65:@7992.4]
  assign _T_8595 = _T_8565[29]; // @[Bitwise.scala 50:65:@7993.4]
  assign _T_8596 = _T_8565[30]; // @[Bitwise.scala 50:65:@7994.4]
  assign _T_8597 = _T_8565[31]; // @[Bitwise.scala 50:65:@7995.4]
  assign _T_8598 = _T_8565[32]; // @[Bitwise.scala 50:65:@7996.4]
  assign _T_8599 = _T_8565[33]; // @[Bitwise.scala 50:65:@7997.4]
  assign _T_8600 = _T_8565[34]; // @[Bitwise.scala 50:65:@7998.4]
  assign _T_8601 = _T_8565[35]; // @[Bitwise.scala 50:65:@7999.4]
  assign _T_8602 = _T_8565[36]; // @[Bitwise.scala 50:65:@8000.4]
  assign _T_8603 = _T_8565[37]; // @[Bitwise.scala 50:65:@8001.4]
  assign _T_8604 = _T_8565[38]; // @[Bitwise.scala 50:65:@8002.4]
  assign _T_8605 = _T_8565[39]; // @[Bitwise.scala 50:65:@8003.4]
  assign _T_8606 = _T_8565[40]; // @[Bitwise.scala 50:65:@8004.4]
  assign _T_8607 = _T_8565[41]; // @[Bitwise.scala 50:65:@8005.4]
  assign _T_8608 = _T_8565[42]; // @[Bitwise.scala 50:65:@8006.4]
  assign _T_8609 = _T_8565[43]; // @[Bitwise.scala 50:65:@8007.4]
  assign _T_8610 = _T_8565[44]; // @[Bitwise.scala 50:65:@8008.4]
  assign _T_8611 = _T_8565[45]; // @[Bitwise.scala 50:65:@8009.4]
  assign _T_8612 = _T_8565[46]; // @[Bitwise.scala 50:65:@8010.4]
  assign _T_8613 = _T_8565[47]; // @[Bitwise.scala 50:65:@8011.4]
  assign _T_8614 = _T_8565[48]; // @[Bitwise.scala 50:65:@8012.4]
  assign _T_8615 = _T_8565[49]; // @[Bitwise.scala 50:65:@8013.4]
  assign _T_8616 = _T_8565[50]; // @[Bitwise.scala 50:65:@8014.4]
  assign _T_8617 = _T_8565[51]; // @[Bitwise.scala 50:65:@8015.4]
  assign _T_8618 = _T_8565[52]; // @[Bitwise.scala 50:65:@8016.4]
  assign _T_8619 = _T_8565[53]; // @[Bitwise.scala 50:65:@8017.4]
  assign _T_8620 = _T_8565[54]; // @[Bitwise.scala 50:65:@8018.4]
  assign _T_8621 = _T_8565[55]; // @[Bitwise.scala 50:65:@8019.4]
  assign _T_8622 = _T_8565[56]; // @[Bitwise.scala 50:65:@8020.4]
  assign _T_8623 = _T_8565[57]; // @[Bitwise.scala 50:65:@8021.4]
  assign _T_8624 = _T_8565[58]; // @[Bitwise.scala 50:65:@8022.4]
  assign _T_8625 = _T_8565[59]; // @[Bitwise.scala 50:65:@8023.4]
  assign _T_8626 = _T_8565[60]; // @[Bitwise.scala 50:65:@8024.4]
  assign _T_8627 = _T_8567 + _T_8568; // @[Bitwise.scala 48:55:@8025.4]
  assign _GEN_991 = {{1'd0}, _T_8566}; // @[Bitwise.scala 48:55:@8026.4]
  assign _T_8628 = _GEN_991 + _T_8627; // @[Bitwise.scala 48:55:@8026.4]
  assign _T_8629 = _T_8569 + _T_8570; // @[Bitwise.scala 48:55:@8027.4]
  assign _T_8630 = _T_8571 + _T_8572; // @[Bitwise.scala 48:55:@8028.4]
  assign _T_8631 = _T_8629 + _T_8630; // @[Bitwise.scala 48:55:@8029.4]
  assign _T_8632 = _T_8628 + _T_8631; // @[Bitwise.scala 48:55:@8030.4]
  assign _T_8633 = _T_8573 + _T_8574; // @[Bitwise.scala 48:55:@8031.4]
  assign _T_8634 = _T_8575 + _T_8576; // @[Bitwise.scala 48:55:@8032.4]
  assign _T_8635 = _T_8633 + _T_8634; // @[Bitwise.scala 48:55:@8033.4]
  assign _T_8636 = _T_8577 + _T_8578; // @[Bitwise.scala 48:55:@8034.4]
  assign _T_8637 = _T_8579 + _T_8580; // @[Bitwise.scala 48:55:@8035.4]
  assign _T_8638 = _T_8636 + _T_8637; // @[Bitwise.scala 48:55:@8036.4]
  assign _T_8639 = _T_8635 + _T_8638; // @[Bitwise.scala 48:55:@8037.4]
  assign _T_8640 = _T_8632 + _T_8639; // @[Bitwise.scala 48:55:@8038.4]
  assign _T_8641 = _T_8582 + _T_8583; // @[Bitwise.scala 48:55:@8039.4]
  assign _GEN_992 = {{1'd0}, _T_8581}; // @[Bitwise.scala 48:55:@8040.4]
  assign _T_8642 = _GEN_992 + _T_8641; // @[Bitwise.scala 48:55:@8040.4]
  assign _T_8643 = _T_8584 + _T_8585; // @[Bitwise.scala 48:55:@8041.4]
  assign _T_8644 = _T_8586 + _T_8587; // @[Bitwise.scala 48:55:@8042.4]
  assign _T_8645 = _T_8643 + _T_8644; // @[Bitwise.scala 48:55:@8043.4]
  assign _T_8646 = _T_8642 + _T_8645; // @[Bitwise.scala 48:55:@8044.4]
  assign _T_8647 = _T_8588 + _T_8589; // @[Bitwise.scala 48:55:@8045.4]
  assign _T_8648 = _T_8590 + _T_8591; // @[Bitwise.scala 48:55:@8046.4]
  assign _T_8649 = _T_8647 + _T_8648; // @[Bitwise.scala 48:55:@8047.4]
  assign _T_8650 = _T_8592 + _T_8593; // @[Bitwise.scala 48:55:@8048.4]
  assign _T_8651 = _T_8594 + _T_8595; // @[Bitwise.scala 48:55:@8049.4]
  assign _T_8652 = _T_8650 + _T_8651; // @[Bitwise.scala 48:55:@8050.4]
  assign _T_8653 = _T_8649 + _T_8652; // @[Bitwise.scala 48:55:@8051.4]
  assign _T_8654 = _T_8646 + _T_8653; // @[Bitwise.scala 48:55:@8052.4]
  assign _T_8655 = _T_8640 + _T_8654; // @[Bitwise.scala 48:55:@8053.4]
  assign _T_8656 = _T_8597 + _T_8598; // @[Bitwise.scala 48:55:@8054.4]
  assign _GEN_993 = {{1'd0}, _T_8596}; // @[Bitwise.scala 48:55:@8055.4]
  assign _T_8657 = _GEN_993 + _T_8656; // @[Bitwise.scala 48:55:@8055.4]
  assign _T_8658 = _T_8599 + _T_8600; // @[Bitwise.scala 48:55:@8056.4]
  assign _T_8659 = _T_8601 + _T_8602; // @[Bitwise.scala 48:55:@8057.4]
  assign _T_8660 = _T_8658 + _T_8659; // @[Bitwise.scala 48:55:@8058.4]
  assign _T_8661 = _T_8657 + _T_8660; // @[Bitwise.scala 48:55:@8059.4]
  assign _T_8662 = _T_8603 + _T_8604; // @[Bitwise.scala 48:55:@8060.4]
  assign _T_8663 = _T_8605 + _T_8606; // @[Bitwise.scala 48:55:@8061.4]
  assign _T_8664 = _T_8662 + _T_8663; // @[Bitwise.scala 48:55:@8062.4]
  assign _T_8665 = _T_8607 + _T_8608; // @[Bitwise.scala 48:55:@8063.4]
  assign _T_8666 = _T_8609 + _T_8610; // @[Bitwise.scala 48:55:@8064.4]
  assign _T_8667 = _T_8665 + _T_8666; // @[Bitwise.scala 48:55:@8065.4]
  assign _T_8668 = _T_8664 + _T_8667; // @[Bitwise.scala 48:55:@8066.4]
  assign _T_8669 = _T_8661 + _T_8668; // @[Bitwise.scala 48:55:@8067.4]
  assign _T_8670 = _T_8611 + _T_8612; // @[Bitwise.scala 48:55:@8068.4]
  assign _T_8671 = _T_8613 + _T_8614; // @[Bitwise.scala 48:55:@8069.4]
  assign _T_8672 = _T_8670 + _T_8671; // @[Bitwise.scala 48:55:@8070.4]
  assign _T_8673 = _T_8615 + _T_8616; // @[Bitwise.scala 48:55:@8071.4]
  assign _T_8674 = _T_8617 + _T_8618; // @[Bitwise.scala 48:55:@8072.4]
  assign _T_8675 = _T_8673 + _T_8674; // @[Bitwise.scala 48:55:@8073.4]
  assign _T_8676 = _T_8672 + _T_8675; // @[Bitwise.scala 48:55:@8074.4]
  assign _T_8677 = _T_8619 + _T_8620; // @[Bitwise.scala 48:55:@8075.4]
  assign _T_8678 = _T_8621 + _T_8622; // @[Bitwise.scala 48:55:@8076.4]
  assign _T_8679 = _T_8677 + _T_8678; // @[Bitwise.scala 48:55:@8077.4]
  assign _T_8680 = _T_8623 + _T_8624; // @[Bitwise.scala 48:55:@8078.4]
  assign _T_8681 = _T_8625 + _T_8626; // @[Bitwise.scala 48:55:@8079.4]
  assign _T_8682 = _T_8680 + _T_8681; // @[Bitwise.scala 48:55:@8080.4]
  assign _T_8683 = _T_8679 + _T_8682; // @[Bitwise.scala 48:55:@8081.4]
  assign _T_8684 = _T_8676 + _T_8683; // @[Bitwise.scala 48:55:@8082.4]
  assign _T_8685 = _T_8669 + _T_8684; // @[Bitwise.scala 48:55:@8083.4]
  assign _T_8686 = _T_8655 + _T_8685; // @[Bitwise.scala 48:55:@8084.4]
  assign _T_8750 = _T_1124[61:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@8149.4]
  assign _T_8751 = _T_8750[0]; // @[Bitwise.scala 50:65:@8150.4]
  assign _T_8752 = _T_8750[1]; // @[Bitwise.scala 50:65:@8151.4]
  assign _T_8753 = _T_8750[2]; // @[Bitwise.scala 50:65:@8152.4]
  assign _T_8754 = _T_8750[3]; // @[Bitwise.scala 50:65:@8153.4]
  assign _T_8755 = _T_8750[4]; // @[Bitwise.scala 50:65:@8154.4]
  assign _T_8756 = _T_8750[5]; // @[Bitwise.scala 50:65:@8155.4]
  assign _T_8757 = _T_8750[6]; // @[Bitwise.scala 50:65:@8156.4]
  assign _T_8758 = _T_8750[7]; // @[Bitwise.scala 50:65:@8157.4]
  assign _T_8759 = _T_8750[8]; // @[Bitwise.scala 50:65:@8158.4]
  assign _T_8760 = _T_8750[9]; // @[Bitwise.scala 50:65:@8159.4]
  assign _T_8761 = _T_8750[10]; // @[Bitwise.scala 50:65:@8160.4]
  assign _T_8762 = _T_8750[11]; // @[Bitwise.scala 50:65:@8161.4]
  assign _T_8763 = _T_8750[12]; // @[Bitwise.scala 50:65:@8162.4]
  assign _T_8764 = _T_8750[13]; // @[Bitwise.scala 50:65:@8163.4]
  assign _T_8765 = _T_8750[14]; // @[Bitwise.scala 50:65:@8164.4]
  assign _T_8766 = _T_8750[15]; // @[Bitwise.scala 50:65:@8165.4]
  assign _T_8767 = _T_8750[16]; // @[Bitwise.scala 50:65:@8166.4]
  assign _T_8768 = _T_8750[17]; // @[Bitwise.scala 50:65:@8167.4]
  assign _T_8769 = _T_8750[18]; // @[Bitwise.scala 50:65:@8168.4]
  assign _T_8770 = _T_8750[19]; // @[Bitwise.scala 50:65:@8169.4]
  assign _T_8771 = _T_8750[20]; // @[Bitwise.scala 50:65:@8170.4]
  assign _T_8772 = _T_8750[21]; // @[Bitwise.scala 50:65:@8171.4]
  assign _T_8773 = _T_8750[22]; // @[Bitwise.scala 50:65:@8172.4]
  assign _T_8774 = _T_8750[23]; // @[Bitwise.scala 50:65:@8173.4]
  assign _T_8775 = _T_8750[24]; // @[Bitwise.scala 50:65:@8174.4]
  assign _T_8776 = _T_8750[25]; // @[Bitwise.scala 50:65:@8175.4]
  assign _T_8777 = _T_8750[26]; // @[Bitwise.scala 50:65:@8176.4]
  assign _T_8778 = _T_8750[27]; // @[Bitwise.scala 50:65:@8177.4]
  assign _T_8779 = _T_8750[28]; // @[Bitwise.scala 50:65:@8178.4]
  assign _T_8780 = _T_8750[29]; // @[Bitwise.scala 50:65:@8179.4]
  assign _T_8781 = _T_8750[30]; // @[Bitwise.scala 50:65:@8180.4]
  assign _T_8782 = _T_8750[31]; // @[Bitwise.scala 50:65:@8181.4]
  assign _T_8783 = _T_8750[32]; // @[Bitwise.scala 50:65:@8182.4]
  assign _T_8784 = _T_8750[33]; // @[Bitwise.scala 50:65:@8183.4]
  assign _T_8785 = _T_8750[34]; // @[Bitwise.scala 50:65:@8184.4]
  assign _T_8786 = _T_8750[35]; // @[Bitwise.scala 50:65:@8185.4]
  assign _T_8787 = _T_8750[36]; // @[Bitwise.scala 50:65:@8186.4]
  assign _T_8788 = _T_8750[37]; // @[Bitwise.scala 50:65:@8187.4]
  assign _T_8789 = _T_8750[38]; // @[Bitwise.scala 50:65:@8188.4]
  assign _T_8790 = _T_8750[39]; // @[Bitwise.scala 50:65:@8189.4]
  assign _T_8791 = _T_8750[40]; // @[Bitwise.scala 50:65:@8190.4]
  assign _T_8792 = _T_8750[41]; // @[Bitwise.scala 50:65:@8191.4]
  assign _T_8793 = _T_8750[42]; // @[Bitwise.scala 50:65:@8192.4]
  assign _T_8794 = _T_8750[43]; // @[Bitwise.scala 50:65:@8193.4]
  assign _T_8795 = _T_8750[44]; // @[Bitwise.scala 50:65:@8194.4]
  assign _T_8796 = _T_8750[45]; // @[Bitwise.scala 50:65:@8195.4]
  assign _T_8797 = _T_8750[46]; // @[Bitwise.scala 50:65:@8196.4]
  assign _T_8798 = _T_8750[47]; // @[Bitwise.scala 50:65:@8197.4]
  assign _T_8799 = _T_8750[48]; // @[Bitwise.scala 50:65:@8198.4]
  assign _T_8800 = _T_8750[49]; // @[Bitwise.scala 50:65:@8199.4]
  assign _T_8801 = _T_8750[50]; // @[Bitwise.scala 50:65:@8200.4]
  assign _T_8802 = _T_8750[51]; // @[Bitwise.scala 50:65:@8201.4]
  assign _T_8803 = _T_8750[52]; // @[Bitwise.scala 50:65:@8202.4]
  assign _T_8804 = _T_8750[53]; // @[Bitwise.scala 50:65:@8203.4]
  assign _T_8805 = _T_8750[54]; // @[Bitwise.scala 50:65:@8204.4]
  assign _T_8806 = _T_8750[55]; // @[Bitwise.scala 50:65:@8205.4]
  assign _T_8807 = _T_8750[56]; // @[Bitwise.scala 50:65:@8206.4]
  assign _T_8808 = _T_8750[57]; // @[Bitwise.scala 50:65:@8207.4]
  assign _T_8809 = _T_8750[58]; // @[Bitwise.scala 50:65:@8208.4]
  assign _T_8810 = _T_8750[59]; // @[Bitwise.scala 50:65:@8209.4]
  assign _T_8811 = _T_8750[60]; // @[Bitwise.scala 50:65:@8210.4]
  assign _T_8812 = _T_8750[61]; // @[Bitwise.scala 50:65:@8211.4]
  assign _T_8813 = _T_8752 + _T_8753; // @[Bitwise.scala 48:55:@8212.4]
  assign _GEN_994 = {{1'd0}, _T_8751}; // @[Bitwise.scala 48:55:@8213.4]
  assign _T_8814 = _GEN_994 + _T_8813; // @[Bitwise.scala 48:55:@8213.4]
  assign _T_8815 = _T_8754 + _T_8755; // @[Bitwise.scala 48:55:@8214.4]
  assign _T_8816 = _T_8756 + _T_8757; // @[Bitwise.scala 48:55:@8215.4]
  assign _T_8817 = _T_8815 + _T_8816; // @[Bitwise.scala 48:55:@8216.4]
  assign _T_8818 = _T_8814 + _T_8817; // @[Bitwise.scala 48:55:@8217.4]
  assign _T_8819 = _T_8758 + _T_8759; // @[Bitwise.scala 48:55:@8218.4]
  assign _T_8820 = _T_8760 + _T_8761; // @[Bitwise.scala 48:55:@8219.4]
  assign _T_8821 = _T_8819 + _T_8820; // @[Bitwise.scala 48:55:@8220.4]
  assign _T_8822 = _T_8762 + _T_8763; // @[Bitwise.scala 48:55:@8221.4]
  assign _T_8823 = _T_8764 + _T_8765; // @[Bitwise.scala 48:55:@8222.4]
  assign _T_8824 = _T_8822 + _T_8823; // @[Bitwise.scala 48:55:@8223.4]
  assign _T_8825 = _T_8821 + _T_8824; // @[Bitwise.scala 48:55:@8224.4]
  assign _T_8826 = _T_8818 + _T_8825; // @[Bitwise.scala 48:55:@8225.4]
  assign _T_8827 = _T_8766 + _T_8767; // @[Bitwise.scala 48:55:@8226.4]
  assign _T_8828 = _T_8768 + _T_8769; // @[Bitwise.scala 48:55:@8227.4]
  assign _T_8829 = _T_8827 + _T_8828; // @[Bitwise.scala 48:55:@8228.4]
  assign _T_8830 = _T_8770 + _T_8771; // @[Bitwise.scala 48:55:@8229.4]
  assign _T_8831 = _T_8772 + _T_8773; // @[Bitwise.scala 48:55:@8230.4]
  assign _T_8832 = _T_8830 + _T_8831; // @[Bitwise.scala 48:55:@8231.4]
  assign _T_8833 = _T_8829 + _T_8832; // @[Bitwise.scala 48:55:@8232.4]
  assign _T_8834 = _T_8774 + _T_8775; // @[Bitwise.scala 48:55:@8233.4]
  assign _T_8835 = _T_8776 + _T_8777; // @[Bitwise.scala 48:55:@8234.4]
  assign _T_8836 = _T_8834 + _T_8835; // @[Bitwise.scala 48:55:@8235.4]
  assign _T_8837 = _T_8778 + _T_8779; // @[Bitwise.scala 48:55:@8236.4]
  assign _T_8838 = _T_8780 + _T_8781; // @[Bitwise.scala 48:55:@8237.4]
  assign _T_8839 = _T_8837 + _T_8838; // @[Bitwise.scala 48:55:@8238.4]
  assign _T_8840 = _T_8836 + _T_8839; // @[Bitwise.scala 48:55:@8239.4]
  assign _T_8841 = _T_8833 + _T_8840; // @[Bitwise.scala 48:55:@8240.4]
  assign _T_8842 = _T_8826 + _T_8841; // @[Bitwise.scala 48:55:@8241.4]
  assign _T_8843 = _T_8783 + _T_8784; // @[Bitwise.scala 48:55:@8242.4]
  assign _GEN_995 = {{1'd0}, _T_8782}; // @[Bitwise.scala 48:55:@8243.4]
  assign _T_8844 = _GEN_995 + _T_8843; // @[Bitwise.scala 48:55:@8243.4]
  assign _T_8845 = _T_8785 + _T_8786; // @[Bitwise.scala 48:55:@8244.4]
  assign _T_8846 = _T_8787 + _T_8788; // @[Bitwise.scala 48:55:@8245.4]
  assign _T_8847 = _T_8845 + _T_8846; // @[Bitwise.scala 48:55:@8246.4]
  assign _T_8848 = _T_8844 + _T_8847; // @[Bitwise.scala 48:55:@8247.4]
  assign _T_8849 = _T_8789 + _T_8790; // @[Bitwise.scala 48:55:@8248.4]
  assign _T_8850 = _T_8791 + _T_8792; // @[Bitwise.scala 48:55:@8249.4]
  assign _T_8851 = _T_8849 + _T_8850; // @[Bitwise.scala 48:55:@8250.4]
  assign _T_8852 = _T_8793 + _T_8794; // @[Bitwise.scala 48:55:@8251.4]
  assign _T_8853 = _T_8795 + _T_8796; // @[Bitwise.scala 48:55:@8252.4]
  assign _T_8854 = _T_8852 + _T_8853; // @[Bitwise.scala 48:55:@8253.4]
  assign _T_8855 = _T_8851 + _T_8854; // @[Bitwise.scala 48:55:@8254.4]
  assign _T_8856 = _T_8848 + _T_8855; // @[Bitwise.scala 48:55:@8255.4]
  assign _T_8857 = _T_8797 + _T_8798; // @[Bitwise.scala 48:55:@8256.4]
  assign _T_8858 = _T_8799 + _T_8800; // @[Bitwise.scala 48:55:@8257.4]
  assign _T_8859 = _T_8857 + _T_8858; // @[Bitwise.scala 48:55:@8258.4]
  assign _T_8860 = _T_8801 + _T_8802; // @[Bitwise.scala 48:55:@8259.4]
  assign _T_8861 = _T_8803 + _T_8804; // @[Bitwise.scala 48:55:@8260.4]
  assign _T_8862 = _T_8860 + _T_8861; // @[Bitwise.scala 48:55:@8261.4]
  assign _T_8863 = _T_8859 + _T_8862; // @[Bitwise.scala 48:55:@8262.4]
  assign _T_8864 = _T_8805 + _T_8806; // @[Bitwise.scala 48:55:@8263.4]
  assign _T_8865 = _T_8807 + _T_8808; // @[Bitwise.scala 48:55:@8264.4]
  assign _T_8866 = _T_8864 + _T_8865; // @[Bitwise.scala 48:55:@8265.4]
  assign _T_8867 = _T_8809 + _T_8810; // @[Bitwise.scala 48:55:@8266.4]
  assign _T_8868 = _T_8811 + _T_8812; // @[Bitwise.scala 48:55:@8267.4]
  assign _T_8869 = _T_8867 + _T_8868; // @[Bitwise.scala 48:55:@8268.4]
  assign _T_8870 = _T_8866 + _T_8869; // @[Bitwise.scala 48:55:@8269.4]
  assign _T_8871 = _T_8863 + _T_8870; // @[Bitwise.scala 48:55:@8270.4]
  assign _T_8872 = _T_8856 + _T_8871; // @[Bitwise.scala 48:55:@8271.4]
  assign _T_8873 = _T_8842 + _T_8872; // @[Bitwise.scala 48:55:@8272.4]
  assign _T_8937 = _T_1124[62:0]; // @[NV_NVDLA_CSC_WL_dec.scala 85:60:@8337.4]
  assign _T_8938 = _T_8937[0]; // @[Bitwise.scala 50:65:@8338.4]
  assign _T_8939 = _T_8937[1]; // @[Bitwise.scala 50:65:@8339.4]
  assign _T_8940 = _T_8937[2]; // @[Bitwise.scala 50:65:@8340.4]
  assign _T_8941 = _T_8937[3]; // @[Bitwise.scala 50:65:@8341.4]
  assign _T_8942 = _T_8937[4]; // @[Bitwise.scala 50:65:@8342.4]
  assign _T_8943 = _T_8937[5]; // @[Bitwise.scala 50:65:@8343.4]
  assign _T_8944 = _T_8937[6]; // @[Bitwise.scala 50:65:@8344.4]
  assign _T_8945 = _T_8937[7]; // @[Bitwise.scala 50:65:@8345.4]
  assign _T_8946 = _T_8937[8]; // @[Bitwise.scala 50:65:@8346.4]
  assign _T_8947 = _T_8937[9]; // @[Bitwise.scala 50:65:@8347.4]
  assign _T_8948 = _T_8937[10]; // @[Bitwise.scala 50:65:@8348.4]
  assign _T_8949 = _T_8937[11]; // @[Bitwise.scala 50:65:@8349.4]
  assign _T_8950 = _T_8937[12]; // @[Bitwise.scala 50:65:@8350.4]
  assign _T_8951 = _T_8937[13]; // @[Bitwise.scala 50:65:@8351.4]
  assign _T_8952 = _T_8937[14]; // @[Bitwise.scala 50:65:@8352.4]
  assign _T_8953 = _T_8937[15]; // @[Bitwise.scala 50:65:@8353.4]
  assign _T_8954 = _T_8937[16]; // @[Bitwise.scala 50:65:@8354.4]
  assign _T_8955 = _T_8937[17]; // @[Bitwise.scala 50:65:@8355.4]
  assign _T_8956 = _T_8937[18]; // @[Bitwise.scala 50:65:@8356.4]
  assign _T_8957 = _T_8937[19]; // @[Bitwise.scala 50:65:@8357.4]
  assign _T_8958 = _T_8937[20]; // @[Bitwise.scala 50:65:@8358.4]
  assign _T_8959 = _T_8937[21]; // @[Bitwise.scala 50:65:@8359.4]
  assign _T_8960 = _T_8937[22]; // @[Bitwise.scala 50:65:@8360.4]
  assign _T_8961 = _T_8937[23]; // @[Bitwise.scala 50:65:@8361.4]
  assign _T_8962 = _T_8937[24]; // @[Bitwise.scala 50:65:@8362.4]
  assign _T_8963 = _T_8937[25]; // @[Bitwise.scala 50:65:@8363.4]
  assign _T_8964 = _T_8937[26]; // @[Bitwise.scala 50:65:@8364.4]
  assign _T_8965 = _T_8937[27]; // @[Bitwise.scala 50:65:@8365.4]
  assign _T_8966 = _T_8937[28]; // @[Bitwise.scala 50:65:@8366.4]
  assign _T_8967 = _T_8937[29]; // @[Bitwise.scala 50:65:@8367.4]
  assign _T_8968 = _T_8937[30]; // @[Bitwise.scala 50:65:@8368.4]
  assign _T_8969 = _T_8937[31]; // @[Bitwise.scala 50:65:@8369.4]
  assign _T_8970 = _T_8937[32]; // @[Bitwise.scala 50:65:@8370.4]
  assign _T_8971 = _T_8937[33]; // @[Bitwise.scala 50:65:@8371.4]
  assign _T_8972 = _T_8937[34]; // @[Bitwise.scala 50:65:@8372.4]
  assign _T_8973 = _T_8937[35]; // @[Bitwise.scala 50:65:@8373.4]
  assign _T_8974 = _T_8937[36]; // @[Bitwise.scala 50:65:@8374.4]
  assign _T_8975 = _T_8937[37]; // @[Bitwise.scala 50:65:@8375.4]
  assign _T_8976 = _T_8937[38]; // @[Bitwise.scala 50:65:@8376.4]
  assign _T_8977 = _T_8937[39]; // @[Bitwise.scala 50:65:@8377.4]
  assign _T_8978 = _T_8937[40]; // @[Bitwise.scala 50:65:@8378.4]
  assign _T_8979 = _T_8937[41]; // @[Bitwise.scala 50:65:@8379.4]
  assign _T_8980 = _T_8937[42]; // @[Bitwise.scala 50:65:@8380.4]
  assign _T_8981 = _T_8937[43]; // @[Bitwise.scala 50:65:@8381.4]
  assign _T_8982 = _T_8937[44]; // @[Bitwise.scala 50:65:@8382.4]
  assign _T_8983 = _T_8937[45]; // @[Bitwise.scala 50:65:@8383.4]
  assign _T_8984 = _T_8937[46]; // @[Bitwise.scala 50:65:@8384.4]
  assign _T_8985 = _T_8937[47]; // @[Bitwise.scala 50:65:@8385.4]
  assign _T_8986 = _T_8937[48]; // @[Bitwise.scala 50:65:@8386.4]
  assign _T_8987 = _T_8937[49]; // @[Bitwise.scala 50:65:@8387.4]
  assign _T_8988 = _T_8937[50]; // @[Bitwise.scala 50:65:@8388.4]
  assign _T_8989 = _T_8937[51]; // @[Bitwise.scala 50:65:@8389.4]
  assign _T_8990 = _T_8937[52]; // @[Bitwise.scala 50:65:@8390.4]
  assign _T_8991 = _T_8937[53]; // @[Bitwise.scala 50:65:@8391.4]
  assign _T_8992 = _T_8937[54]; // @[Bitwise.scala 50:65:@8392.4]
  assign _T_8993 = _T_8937[55]; // @[Bitwise.scala 50:65:@8393.4]
  assign _T_8994 = _T_8937[56]; // @[Bitwise.scala 50:65:@8394.4]
  assign _T_8995 = _T_8937[57]; // @[Bitwise.scala 50:65:@8395.4]
  assign _T_8996 = _T_8937[58]; // @[Bitwise.scala 50:65:@8396.4]
  assign _T_8997 = _T_8937[59]; // @[Bitwise.scala 50:65:@8397.4]
  assign _T_8998 = _T_8937[60]; // @[Bitwise.scala 50:65:@8398.4]
  assign _T_8999 = _T_8937[61]; // @[Bitwise.scala 50:65:@8399.4]
  assign _T_9000 = _T_8937[62]; // @[Bitwise.scala 50:65:@8400.4]
  assign _T_9001 = _T_8939 + _T_8940; // @[Bitwise.scala 48:55:@8401.4]
  assign _GEN_996 = {{1'd0}, _T_8938}; // @[Bitwise.scala 48:55:@8402.4]
  assign _T_9002 = _GEN_996 + _T_9001; // @[Bitwise.scala 48:55:@8402.4]
  assign _T_9003 = _T_8941 + _T_8942; // @[Bitwise.scala 48:55:@8403.4]
  assign _T_9004 = _T_8943 + _T_8944; // @[Bitwise.scala 48:55:@8404.4]
  assign _T_9005 = _T_9003 + _T_9004; // @[Bitwise.scala 48:55:@8405.4]
  assign _T_9006 = _T_9002 + _T_9005; // @[Bitwise.scala 48:55:@8406.4]
  assign _T_9007 = _T_8945 + _T_8946; // @[Bitwise.scala 48:55:@8407.4]
  assign _T_9008 = _T_8947 + _T_8948; // @[Bitwise.scala 48:55:@8408.4]
  assign _T_9009 = _T_9007 + _T_9008; // @[Bitwise.scala 48:55:@8409.4]
  assign _T_9010 = _T_8949 + _T_8950; // @[Bitwise.scala 48:55:@8410.4]
  assign _T_9011 = _T_8951 + _T_8952; // @[Bitwise.scala 48:55:@8411.4]
  assign _T_9012 = _T_9010 + _T_9011; // @[Bitwise.scala 48:55:@8412.4]
  assign _T_9013 = _T_9009 + _T_9012; // @[Bitwise.scala 48:55:@8413.4]
  assign _T_9014 = _T_9006 + _T_9013; // @[Bitwise.scala 48:55:@8414.4]
  assign _T_9015 = _T_8953 + _T_8954; // @[Bitwise.scala 48:55:@8415.4]
  assign _T_9016 = _T_8955 + _T_8956; // @[Bitwise.scala 48:55:@8416.4]
  assign _T_9017 = _T_9015 + _T_9016; // @[Bitwise.scala 48:55:@8417.4]
  assign _T_9018 = _T_8957 + _T_8958; // @[Bitwise.scala 48:55:@8418.4]
  assign _T_9019 = _T_8959 + _T_8960; // @[Bitwise.scala 48:55:@8419.4]
  assign _T_9020 = _T_9018 + _T_9019; // @[Bitwise.scala 48:55:@8420.4]
  assign _T_9021 = _T_9017 + _T_9020; // @[Bitwise.scala 48:55:@8421.4]
  assign _T_9022 = _T_8961 + _T_8962; // @[Bitwise.scala 48:55:@8422.4]
  assign _T_9023 = _T_8963 + _T_8964; // @[Bitwise.scala 48:55:@8423.4]
  assign _T_9024 = _T_9022 + _T_9023; // @[Bitwise.scala 48:55:@8424.4]
  assign _T_9025 = _T_8965 + _T_8966; // @[Bitwise.scala 48:55:@8425.4]
  assign _T_9026 = _T_8967 + _T_8968; // @[Bitwise.scala 48:55:@8426.4]
  assign _T_9027 = _T_9025 + _T_9026; // @[Bitwise.scala 48:55:@8427.4]
  assign _T_9028 = _T_9024 + _T_9027; // @[Bitwise.scala 48:55:@8428.4]
  assign _T_9029 = _T_9021 + _T_9028; // @[Bitwise.scala 48:55:@8429.4]
  assign _T_9030 = _T_9014 + _T_9029; // @[Bitwise.scala 48:55:@8430.4]
  assign _T_9031 = _T_8969 + _T_8970; // @[Bitwise.scala 48:55:@8431.4]
  assign _T_9032 = _T_8971 + _T_8972; // @[Bitwise.scala 48:55:@8432.4]
  assign _T_9033 = _T_9031 + _T_9032; // @[Bitwise.scala 48:55:@8433.4]
  assign _T_9034 = _T_8973 + _T_8974; // @[Bitwise.scala 48:55:@8434.4]
  assign _T_9035 = _T_8975 + _T_8976; // @[Bitwise.scala 48:55:@8435.4]
  assign _T_9036 = _T_9034 + _T_9035; // @[Bitwise.scala 48:55:@8436.4]
  assign _T_9037 = _T_9033 + _T_9036; // @[Bitwise.scala 48:55:@8437.4]
  assign _T_9038 = _T_8977 + _T_8978; // @[Bitwise.scala 48:55:@8438.4]
  assign _T_9039 = _T_8979 + _T_8980; // @[Bitwise.scala 48:55:@8439.4]
  assign _T_9040 = _T_9038 + _T_9039; // @[Bitwise.scala 48:55:@8440.4]
  assign _T_9041 = _T_8981 + _T_8982; // @[Bitwise.scala 48:55:@8441.4]
  assign _T_9042 = _T_8983 + _T_8984; // @[Bitwise.scala 48:55:@8442.4]
  assign _T_9043 = _T_9041 + _T_9042; // @[Bitwise.scala 48:55:@8443.4]
  assign _T_9044 = _T_9040 + _T_9043; // @[Bitwise.scala 48:55:@8444.4]
  assign _T_9045 = _T_9037 + _T_9044; // @[Bitwise.scala 48:55:@8445.4]
  assign _T_9046 = _T_8985 + _T_8986; // @[Bitwise.scala 48:55:@8446.4]
  assign _T_9047 = _T_8987 + _T_8988; // @[Bitwise.scala 48:55:@8447.4]
  assign _T_9048 = _T_9046 + _T_9047; // @[Bitwise.scala 48:55:@8448.4]
  assign _T_9049 = _T_8989 + _T_8990; // @[Bitwise.scala 48:55:@8449.4]
  assign _T_9050 = _T_8991 + _T_8992; // @[Bitwise.scala 48:55:@8450.4]
  assign _T_9051 = _T_9049 + _T_9050; // @[Bitwise.scala 48:55:@8451.4]
  assign _T_9052 = _T_9048 + _T_9051; // @[Bitwise.scala 48:55:@8452.4]
  assign _T_9053 = _T_8993 + _T_8994; // @[Bitwise.scala 48:55:@8453.4]
  assign _T_9054 = _T_8995 + _T_8996; // @[Bitwise.scala 48:55:@8454.4]
  assign _T_9055 = _T_9053 + _T_9054; // @[Bitwise.scala 48:55:@8455.4]
  assign _T_9056 = _T_8997 + _T_8998; // @[Bitwise.scala 48:55:@8456.4]
  assign _T_9057 = _T_8999 + _T_9000; // @[Bitwise.scala 48:55:@8457.4]
  assign _T_9058 = _T_9056 + _T_9057; // @[Bitwise.scala 48:55:@8458.4]
  assign _T_9059 = _T_9055 + _T_9058; // @[Bitwise.scala 48:55:@8459.4]
  assign _T_9060 = _T_9052 + _T_9059; // @[Bitwise.scala 48:55:@8460.4]
  assign _T_9061 = _T_9045 + _T_9060; // @[Bitwise.scala 48:55:@8461.4]
  assign _T_9062 = _T_9030 + _T_9061; // @[Bitwise.scala 48:55:@8462.4]
  assign _T_9128 = _T_1124[1]; // @[Bitwise.scala 50:65:@8529.4]
  assign _T_9129 = _T_1124[2]; // @[Bitwise.scala 50:65:@8530.4]
  assign _T_9130 = _T_1124[3]; // @[Bitwise.scala 50:65:@8531.4]
  assign _T_9131 = _T_1124[4]; // @[Bitwise.scala 50:65:@8532.4]
  assign _T_9132 = _T_1124[5]; // @[Bitwise.scala 50:65:@8533.4]
  assign _T_9133 = _T_1124[6]; // @[Bitwise.scala 50:65:@8534.4]
  assign _T_9134 = _T_1124[7]; // @[Bitwise.scala 50:65:@8535.4]
  assign _T_9135 = _T_1124[8]; // @[Bitwise.scala 50:65:@8536.4]
  assign _T_9136 = _T_1124[9]; // @[Bitwise.scala 50:65:@8537.4]
  assign _T_9137 = _T_1124[10]; // @[Bitwise.scala 50:65:@8538.4]
  assign _T_9138 = _T_1124[11]; // @[Bitwise.scala 50:65:@8539.4]
  assign _T_9139 = _T_1124[12]; // @[Bitwise.scala 50:65:@8540.4]
  assign _T_9140 = _T_1124[13]; // @[Bitwise.scala 50:65:@8541.4]
  assign _T_9141 = _T_1124[14]; // @[Bitwise.scala 50:65:@8542.4]
  assign _T_9142 = _T_1124[15]; // @[Bitwise.scala 50:65:@8543.4]
  assign _T_9143 = _T_1124[16]; // @[Bitwise.scala 50:65:@8544.4]
  assign _T_9144 = _T_1124[17]; // @[Bitwise.scala 50:65:@8545.4]
  assign _T_9145 = _T_1124[18]; // @[Bitwise.scala 50:65:@8546.4]
  assign _T_9146 = _T_1124[19]; // @[Bitwise.scala 50:65:@8547.4]
  assign _T_9147 = _T_1124[20]; // @[Bitwise.scala 50:65:@8548.4]
  assign _T_9148 = _T_1124[21]; // @[Bitwise.scala 50:65:@8549.4]
  assign _T_9149 = _T_1124[22]; // @[Bitwise.scala 50:65:@8550.4]
  assign _T_9150 = _T_1124[23]; // @[Bitwise.scala 50:65:@8551.4]
  assign _T_9151 = _T_1124[24]; // @[Bitwise.scala 50:65:@8552.4]
  assign _T_9152 = _T_1124[25]; // @[Bitwise.scala 50:65:@8553.4]
  assign _T_9153 = _T_1124[26]; // @[Bitwise.scala 50:65:@8554.4]
  assign _T_9154 = _T_1124[27]; // @[Bitwise.scala 50:65:@8555.4]
  assign _T_9155 = _T_1124[28]; // @[Bitwise.scala 50:65:@8556.4]
  assign _T_9156 = _T_1124[29]; // @[Bitwise.scala 50:65:@8557.4]
  assign _T_9157 = _T_1124[30]; // @[Bitwise.scala 50:65:@8558.4]
  assign _T_9158 = _T_1124[31]; // @[Bitwise.scala 50:65:@8559.4]
  assign _T_9159 = _T_1124[32]; // @[Bitwise.scala 50:65:@8560.4]
  assign _T_9160 = _T_1124[33]; // @[Bitwise.scala 50:65:@8561.4]
  assign _T_9161 = _T_1124[34]; // @[Bitwise.scala 50:65:@8562.4]
  assign _T_9162 = _T_1124[35]; // @[Bitwise.scala 50:65:@8563.4]
  assign _T_9163 = _T_1124[36]; // @[Bitwise.scala 50:65:@8564.4]
  assign _T_9164 = _T_1124[37]; // @[Bitwise.scala 50:65:@8565.4]
  assign _T_9165 = _T_1124[38]; // @[Bitwise.scala 50:65:@8566.4]
  assign _T_9166 = _T_1124[39]; // @[Bitwise.scala 50:65:@8567.4]
  assign _T_9167 = _T_1124[40]; // @[Bitwise.scala 50:65:@8568.4]
  assign _T_9168 = _T_1124[41]; // @[Bitwise.scala 50:65:@8569.4]
  assign _T_9169 = _T_1124[42]; // @[Bitwise.scala 50:65:@8570.4]
  assign _T_9170 = _T_1124[43]; // @[Bitwise.scala 50:65:@8571.4]
  assign _T_9171 = _T_1124[44]; // @[Bitwise.scala 50:65:@8572.4]
  assign _T_9172 = _T_1124[45]; // @[Bitwise.scala 50:65:@8573.4]
  assign _T_9173 = _T_1124[46]; // @[Bitwise.scala 50:65:@8574.4]
  assign _T_9174 = _T_1124[47]; // @[Bitwise.scala 50:65:@8575.4]
  assign _T_9175 = _T_1124[48]; // @[Bitwise.scala 50:65:@8576.4]
  assign _T_9176 = _T_1124[49]; // @[Bitwise.scala 50:65:@8577.4]
  assign _T_9177 = _T_1124[50]; // @[Bitwise.scala 50:65:@8578.4]
  assign _T_9178 = _T_1124[51]; // @[Bitwise.scala 50:65:@8579.4]
  assign _T_9179 = _T_1124[52]; // @[Bitwise.scala 50:65:@8580.4]
  assign _T_9180 = _T_1124[53]; // @[Bitwise.scala 50:65:@8581.4]
  assign _T_9181 = _T_1124[54]; // @[Bitwise.scala 50:65:@8582.4]
  assign _T_9182 = _T_1124[55]; // @[Bitwise.scala 50:65:@8583.4]
  assign _T_9183 = _T_1124[56]; // @[Bitwise.scala 50:65:@8584.4]
  assign _T_9184 = _T_1124[57]; // @[Bitwise.scala 50:65:@8585.4]
  assign _T_9185 = _T_1124[58]; // @[Bitwise.scala 50:65:@8586.4]
  assign _T_9186 = _T_1124[59]; // @[Bitwise.scala 50:65:@8587.4]
  assign _T_9187 = _T_1124[60]; // @[Bitwise.scala 50:65:@8588.4]
  assign _T_9188 = _T_1124[61]; // @[Bitwise.scala 50:65:@8589.4]
  assign _T_9189 = _T_1124[62]; // @[Bitwise.scala 50:65:@8590.4]
  assign _T_9190 = _T_1124[63]; // @[Bitwise.scala 50:65:@8591.4]
  assign _T_9191 = _T_1125 + _T_9128; // @[Bitwise.scala 48:55:@8592.4]
  assign _T_9192 = _T_9129 + _T_9130; // @[Bitwise.scala 48:55:@8593.4]
  assign _T_9193 = _T_9191 + _T_9192; // @[Bitwise.scala 48:55:@8594.4]
  assign _T_9194 = _T_9131 + _T_9132; // @[Bitwise.scala 48:55:@8595.4]
  assign _T_9195 = _T_9133 + _T_9134; // @[Bitwise.scala 48:55:@8596.4]
  assign _T_9196 = _T_9194 + _T_9195; // @[Bitwise.scala 48:55:@8597.4]
  assign _T_9197 = _T_9193 + _T_9196; // @[Bitwise.scala 48:55:@8598.4]
  assign _T_9198 = _T_9135 + _T_9136; // @[Bitwise.scala 48:55:@8599.4]
  assign _T_9199 = _T_9137 + _T_9138; // @[Bitwise.scala 48:55:@8600.4]
  assign _T_9200 = _T_9198 + _T_9199; // @[Bitwise.scala 48:55:@8601.4]
  assign _T_9201 = _T_9139 + _T_9140; // @[Bitwise.scala 48:55:@8602.4]
  assign _T_9202 = _T_9141 + _T_9142; // @[Bitwise.scala 48:55:@8603.4]
  assign _T_9203 = _T_9201 + _T_9202; // @[Bitwise.scala 48:55:@8604.4]
  assign _T_9204 = _T_9200 + _T_9203; // @[Bitwise.scala 48:55:@8605.4]
  assign _T_9205 = _T_9197 + _T_9204; // @[Bitwise.scala 48:55:@8606.4]
  assign _T_9206 = _T_9143 + _T_9144; // @[Bitwise.scala 48:55:@8607.4]
  assign _T_9207 = _T_9145 + _T_9146; // @[Bitwise.scala 48:55:@8608.4]
  assign _T_9208 = _T_9206 + _T_9207; // @[Bitwise.scala 48:55:@8609.4]
  assign _T_9209 = _T_9147 + _T_9148; // @[Bitwise.scala 48:55:@8610.4]
  assign _T_9210 = _T_9149 + _T_9150; // @[Bitwise.scala 48:55:@8611.4]
  assign _T_9211 = _T_9209 + _T_9210; // @[Bitwise.scala 48:55:@8612.4]
  assign _T_9212 = _T_9208 + _T_9211; // @[Bitwise.scala 48:55:@8613.4]
  assign _T_9213 = _T_9151 + _T_9152; // @[Bitwise.scala 48:55:@8614.4]
  assign _T_9214 = _T_9153 + _T_9154; // @[Bitwise.scala 48:55:@8615.4]
  assign _T_9215 = _T_9213 + _T_9214; // @[Bitwise.scala 48:55:@8616.4]
  assign _T_9216 = _T_9155 + _T_9156; // @[Bitwise.scala 48:55:@8617.4]
  assign _T_9217 = _T_9157 + _T_9158; // @[Bitwise.scala 48:55:@8618.4]
  assign _T_9218 = _T_9216 + _T_9217; // @[Bitwise.scala 48:55:@8619.4]
  assign _T_9219 = _T_9215 + _T_9218; // @[Bitwise.scala 48:55:@8620.4]
  assign _T_9220 = _T_9212 + _T_9219; // @[Bitwise.scala 48:55:@8621.4]
  assign _T_9221 = _T_9205 + _T_9220; // @[Bitwise.scala 48:55:@8622.4]
  assign _T_9222 = _T_9159 + _T_9160; // @[Bitwise.scala 48:55:@8623.4]
  assign _T_9223 = _T_9161 + _T_9162; // @[Bitwise.scala 48:55:@8624.4]
  assign _T_9224 = _T_9222 + _T_9223; // @[Bitwise.scala 48:55:@8625.4]
  assign _T_9225 = _T_9163 + _T_9164; // @[Bitwise.scala 48:55:@8626.4]
  assign _T_9226 = _T_9165 + _T_9166; // @[Bitwise.scala 48:55:@8627.4]
  assign _T_9227 = _T_9225 + _T_9226; // @[Bitwise.scala 48:55:@8628.4]
  assign _T_9228 = _T_9224 + _T_9227; // @[Bitwise.scala 48:55:@8629.4]
  assign _T_9229 = _T_9167 + _T_9168; // @[Bitwise.scala 48:55:@8630.4]
  assign _T_9230 = _T_9169 + _T_9170; // @[Bitwise.scala 48:55:@8631.4]
  assign _T_9231 = _T_9229 + _T_9230; // @[Bitwise.scala 48:55:@8632.4]
  assign _T_9232 = _T_9171 + _T_9172; // @[Bitwise.scala 48:55:@8633.4]
  assign _T_9233 = _T_9173 + _T_9174; // @[Bitwise.scala 48:55:@8634.4]
  assign _T_9234 = _T_9232 + _T_9233; // @[Bitwise.scala 48:55:@8635.4]
  assign _T_9235 = _T_9231 + _T_9234; // @[Bitwise.scala 48:55:@8636.4]
  assign _T_9236 = _T_9228 + _T_9235; // @[Bitwise.scala 48:55:@8637.4]
  assign _T_9237 = _T_9175 + _T_9176; // @[Bitwise.scala 48:55:@8638.4]
  assign _T_9238 = _T_9177 + _T_9178; // @[Bitwise.scala 48:55:@8639.4]
  assign _T_9239 = _T_9237 + _T_9238; // @[Bitwise.scala 48:55:@8640.4]
  assign _T_9240 = _T_9179 + _T_9180; // @[Bitwise.scala 48:55:@8641.4]
  assign _T_9241 = _T_9181 + _T_9182; // @[Bitwise.scala 48:55:@8642.4]
  assign _T_9242 = _T_9240 + _T_9241; // @[Bitwise.scala 48:55:@8643.4]
  assign _T_9243 = _T_9239 + _T_9242; // @[Bitwise.scala 48:55:@8644.4]
  assign _T_9244 = _T_9183 + _T_9184; // @[Bitwise.scala 48:55:@8645.4]
  assign _T_9245 = _T_9185 + _T_9186; // @[Bitwise.scala 48:55:@8646.4]
  assign _T_9246 = _T_9244 + _T_9245; // @[Bitwise.scala 48:55:@8647.4]
  assign _T_9247 = _T_9187 + _T_9188; // @[Bitwise.scala 48:55:@8648.4]
  assign _T_9248 = _T_9189 + _T_9190; // @[Bitwise.scala 48:55:@8649.4]
  assign _T_9249 = _T_9247 + _T_9248; // @[Bitwise.scala 48:55:@8650.4]
  assign _T_9250 = _T_9246 + _T_9249; // @[Bitwise.scala 48:55:@8651.4]
  assign _T_9251 = _T_9243 + _T_9250; // @[Bitwise.scala 48:55:@8652.4]
  assign _T_9252 = _T_9236 + _T_9251; // @[Bitwise.scala 48:55:@8653.4]
  assign _T_9253 = _T_9221 + _T_9252; // @[Bitwise.scala 48:55:@8654.4]
  assign _GEN_128 = io_input_valid ? _T_633 : _T_9535_0; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_129 = io_input_valid ? _T_634 : _T_9535_1; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_130 = io_input_valid ? _T_635 : _T_9535_2; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_131 = io_input_valid ? _T_636 : _T_9535_3; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_132 = io_input_valid ? _T_637 : _T_9535_4; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_133 = io_input_valid ? _T_638 : _T_9535_5; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_134 = io_input_valid ? _T_639 : _T_9535_6; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_135 = io_input_valid ? _T_640 : _T_9535_7; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_136 = io_input_valid ? _T_641 : _T_9535_8; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_137 = io_input_valid ? _T_642 : _T_9535_9; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_138 = io_input_valid ? _T_643 : _T_9535_10; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_139 = io_input_valid ? _T_644 : _T_9535_11; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_140 = io_input_valid ? _T_645 : _T_9535_12; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_141 = io_input_valid ? _T_646 : _T_9535_13; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_142 = io_input_valid ? _T_647 : _T_9535_14; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_143 = io_input_valid ? _T_648 : _T_9535_15; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_144 = io_input_valid ? _T_649 : _T_9535_16; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_145 = io_input_valid ? _T_650 : _T_9535_17; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_146 = io_input_valid ? _T_651 : _T_9535_18; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_147 = io_input_valid ? _T_652 : _T_9535_19; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_148 = io_input_valid ? _T_653 : _T_9535_20; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_149 = io_input_valid ? _T_654 : _T_9535_21; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_150 = io_input_valid ? _T_655 : _T_9535_22; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_151 = io_input_valid ? _T_656 : _T_9535_23; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_152 = io_input_valid ? _T_657 : _T_9535_24; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_153 = io_input_valid ? _T_658 : _T_9535_25; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_154 = io_input_valid ? _T_659 : _T_9535_26; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_155 = io_input_valid ? _T_660 : _T_9535_27; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_156 = io_input_valid ? _T_661 : _T_9535_28; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_157 = io_input_valid ? _T_662 : _T_9535_29; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_158 = io_input_valid ? _T_663 : _T_9535_30; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _GEN_159 = io_input_valid ? _T_664 : _T_9535_31; // @[NV_NVDLA_CSC_WL_dec.scala 96:25:@8823.4]
  assign _T_10212 = io_input_mask_en[0]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@8985.4]
  assign _T_10213 = io_input_valid & _T_10212; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@8986.4]
  assign _GEN_160 = _T_10213 ? _T_1125 : _T_10211_0; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@8987.4]
  assign _GEN_161 = _T_10213 ? _T_1193 : _T_10211_1; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@8992.4]
  assign _T_1061_2 = _T_1262[1:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@603.4]
  assign _GEN_162 = _T_10213 ? _T_1061_2 : _T_10211_2; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@8997.4]
  assign _GEN_163 = _T_10213 ? _T_1333 : _T_10211_3; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9002.4]
  assign _T_1061_4 = _T_1406[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@749.4]
  assign _GEN_164 = _T_10213 ? _T_1061_4 : _T_10211_4; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9007.4]
  assign _T_1061_5 = _T_1481[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@825.4]
  assign _GEN_165 = _T_10213 ? _T_1061_5 : _T_10211_5; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9012.4]
  assign _T_1061_6 = _T_1558[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@903.4]
  assign _GEN_166 = _T_10213 ? _T_1061_6 : _T_10211_6; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9017.4]
  assign _GEN_167 = _T_10213 ? _T_1637 : _T_10211_7; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9022.4]
  assign _T_10228 = io_input_mask_en[1]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9025.4]
  assign _T_10229 = io_input_valid & _T_10228; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9026.4]
  assign _T_1061_8 = _T_1718[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1065.4]
  assign _GEN_168 = _T_10229 ? _T_1061_8 : _T_10211_8; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9027.4]
  assign _T_1061_9 = _T_1801[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1149.4]
  assign _GEN_169 = _T_10229 ? _T_1061_9 : _T_10211_9; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9032.4]
  assign _T_1061_10 = _T_1886[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1235.4]
  assign _GEN_170 = _T_10229 ? _T_1061_10 : _T_10211_10; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9037.4]
  assign _T_1061_11 = _T_1973[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1323.4]
  assign _GEN_171 = _T_10229 ? _T_1061_11 : _T_10211_11; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9042.4]
  assign _T_1061_12 = _T_2062[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1413.4]
  assign _GEN_172 = _T_10229 ? _T_1061_12 : _T_10211_12; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9047.4]
  assign _T_1061_13 = _T_2153[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1505.4]
  assign _GEN_173 = _T_10229 ? _T_1061_13 : _T_10211_13; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9052.4]
  assign _T_1061_14 = _T_2246[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1599.4]
  assign _GEN_174 = _T_10229 ? _T_1061_14 : _T_10211_14; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9057.4]
  assign _GEN_175 = _T_10229 ? _T_2341 : _T_10211_15; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9062.4]
  assign _T_10244 = io_input_mask_en[2]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9065.4]
  assign _T_10245 = io_input_valid & _T_10244; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9066.4]
  assign _T_1061_16 = _T_2438[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1793.4]
  assign _GEN_176 = _T_10245 ? _T_1061_16 : _T_10211_16; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9067.4]
  assign _T_1061_17 = _T_2537[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1893.4]
  assign _GEN_177 = _T_10245 ? _T_1061_17 : _T_10211_17; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9072.4]
  assign _T_1061_18 = _T_2638[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@1995.4]
  assign _GEN_178 = _T_10245 ? _T_1061_18 : _T_10211_18; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9077.4]
  assign _T_1061_19 = _T_2741[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2099.4]
  assign _GEN_179 = _T_10245 ? _T_1061_19 : _T_10211_19; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9082.4]
  assign _T_1061_20 = _T_2846[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2205.4]
  assign _GEN_180 = _T_10245 ? _T_1061_20 : _T_10211_20; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9087.4]
  assign _T_1061_21 = _T_2953[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2313.4]
  assign _GEN_181 = _T_10245 ? _T_1061_21 : _T_10211_21; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9092.4]
  assign _T_1061_22 = _T_3062[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2423.4]
  assign _GEN_182 = _T_10245 ? _T_1061_22 : _T_10211_22; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9097.4]
  assign _T_1061_23 = _T_3173[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2535.4]
  assign _GEN_183 = _T_10245 ? _T_1061_23 : _T_10211_23; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9102.4]
  assign _T_10260 = io_input_mask_en[3]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9105.4]
  assign _T_10261 = io_input_valid & _T_10260; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9106.4]
  assign _T_1061_24 = _T_3286[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2649.4]
  assign _GEN_184 = _T_10261 ? _T_1061_24 : _T_10211_24; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9107.4]
  assign _T_1061_25 = _T_3401[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2765.4]
  assign _GEN_185 = _T_10261 ? _T_1061_25 : _T_10211_25; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9112.4]
  assign _T_1061_26 = _T_3518[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@2883.4]
  assign _GEN_186 = _T_10261 ? _T_1061_26 : _T_10211_26; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9117.4]
  assign _T_1061_27 = _T_3637[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3003.4]
  assign _GEN_187 = _T_10261 ? _T_1061_27 : _T_10211_27; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9122.4]
  assign _T_1061_28 = _T_3758[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3125.4]
  assign _GEN_188 = _T_10261 ? _T_1061_28 : _T_10211_28; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9127.4]
  assign _T_1061_29 = _T_3881[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3249.4]
  assign _GEN_189 = _T_10261 ? _T_1061_29 : _T_10211_29; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9132.4]
  assign _T_1061_30 = _T_4006[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3375.4]
  assign _GEN_190 = _T_10261 ? _T_1061_30 : _T_10211_30; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9137.4]
  assign _GEN_191 = _T_10261 ? _T_4133 : _T_10211_31; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9142.4]
  assign _T_10276 = io_input_mask_en[4]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9145.4]
  assign _T_10277 = io_input_valid & _T_10276; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9146.4]
  assign _T_1061_32 = _T_4262[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3633.4]
  assign _GEN_192 = _T_10277 ? _T_1061_32 : _T_10211_32; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9147.4]
  assign _T_1061_33 = _T_4393[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3765.4]
  assign _GEN_193 = _T_10277 ? _T_1061_33 : _T_10211_33; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9152.4]
  assign _T_1061_34 = _T_4526[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@3899.4]
  assign _GEN_194 = _T_10277 ? _T_1061_34 : _T_10211_34; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9157.4]
  assign _T_1061_35 = _T_4661[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4035.4]
  assign _GEN_195 = _T_10277 ? _T_1061_35 : _T_10211_35; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9162.4]
  assign _T_1061_36 = _T_4798[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4173.4]
  assign _GEN_196 = _T_10277 ? _T_1061_36 : _T_10211_36; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9167.4]
  assign _T_1061_37 = _T_4937[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4313.4]
  assign _GEN_197 = _T_10277 ? _T_1061_37 : _T_10211_37; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9172.4]
  assign _T_1061_38 = _T_5078[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4455.4]
  assign _GEN_198 = _T_10277 ? _T_1061_38 : _T_10211_38; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9177.4]
  assign _T_1061_39 = _T_5221[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4599.4]
  assign _GEN_199 = _T_10277 ? _T_1061_39 : _T_10211_39; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9182.4]
  assign _T_10292 = io_input_mask_en[5]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9185.4]
  assign _T_10293 = io_input_valid & _T_10292; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9186.4]
  assign _T_1061_40 = _T_5366[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4745.4]
  assign _GEN_200 = _T_10293 ? _T_1061_40 : _T_10211_40; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9187.4]
  assign _T_1061_41 = _T_5513[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@4893.4]
  assign _GEN_201 = _T_10293 ? _T_1061_41 : _T_10211_41; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9192.4]
  assign _T_1061_42 = _T_5662[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5043.4]
  assign _GEN_202 = _T_10293 ? _T_1061_42 : _T_10211_42; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9197.4]
  assign _T_1061_43 = _T_5813[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5195.4]
  assign _GEN_203 = _T_10293 ? _T_1061_43 : _T_10211_43; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9202.4]
  assign _T_1061_44 = _T_5966[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5349.4]
  assign _GEN_204 = _T_10293 ? _T_1061_44 : _T_10211_44; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9207.4]
  assign _T_1061_45 = _T_6121[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5505.4]
  assign _GEN_205 = _T_10293 ? _T_1061_45 : _T_10211_45; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9212.4]
  assign _T_1061_46 = _T_6278[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5663.4]
  assign _GEN_206 = _T_10293 ? _T_1061_46 : _T_10211_46; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9217.4]
  assign _T_1061_47 = _T_6437[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5823.4]
  assign _GEN_207 = _T_10293 ? _T_1061_47 : _T_10211_47; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9222.4]
  assign _T_10308 = io_input_mask_en[6]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9225.4]
  assign _T_10309 = io_input_valid & _T_10308; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9226.4]
  assign _T_1061_48 = _T_6598[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@5985.4]
  assign _GEN_208 = _T_10309 ? _T_1061_48 : _T_10211_48; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9227.4]
  assign _T_1061_49 = _T_6761[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6149.4]
  assign _GEN_209 = _T_10309 ? _T_1061_49 : _T_10211_49; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9232.4]
  assign _T_1061_50 = _T_6926[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6315.4]
  assign _GEN_210 = _T_10309 ? _T_1061_50 : _T_10211_50; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9237.4]
  assign _T_1061_51 = _T_7093[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6483.4]
  assign _GEN_211 = _T_10309 ? _T_1061_51 : _T_10211_51; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9242.4]
  assign _T_1061_52 = _T_7262[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6653.4]
  assign _GEN_212 = _T_10309 ? _T_1061_52 : _T_10211_52; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9247.4]
  assign _T_1061_53 = _T_7433[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6825.4]
  assign _GEN_213 = _T_10309 ? _T_1061_53 : _T_10211_53; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9252.4]
  assign _T_1061_54 = _T_7606[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@6999.4]
  assign _GEN_214 = _T_10309 ? _T_1061_54 : _T_10211_54; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9257.4]
  assign _T_1061_55 = _T_7781[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7175.4]
  assign _GEN_215 = _T_10309 ? _T_1061_55 : _T_10211_55; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9262.4]
  assign _T_10324 = io_input_mask_en[7]; // @[NV_NVDLA_CSC_WL_dec.scala 103:47:@9265.4]
  assign _T_10325 = io_input_valid & _T_10324; // @[NV_NVDLA_CSC_WL_dec.scala 103:29:@9266.4]
  assign _T_1061_56 = _T_7958[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7353.4]
  assign _GEN_216 = _T_10325 ? _T_1061_56 : _T_10211_56; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9267.4]
  assign _T_1061_57 = _T_8137[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7533.4]
  assign _GEN_217 = _T_10325 ? _T_1061_57 : _T_10211_57; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9272.4]
  assign _T_1061_58 = _T_8318[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7715.4]
  assign _GEN_218 = _T_10325 ? _T_1061_58 : _T_10211_58; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9277.4]
  assign _T_1061_59 = _T_8501[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@7899.4]
  assign _GEN_219 = _T_10325 ? _T_1061_59 : _T_10211_59; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9282.4]
  assign _T_1061_60 = _T_8686[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@8085.4]
  assign _GEN_220 = _T_10325 ? _T_1061_60 : _T_10211_60; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9287.4]
  assign _T_1061_61 = _T_8873[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@8273.4]
  assign _GEN_221 = _T_10325 ? _T_1061_61 : _T_10211_61; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9292.4]
  assign _T_1061_62 = _T_9062[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 82:23:@399.4 NV_NVDLA_CSC_WL_dec.scala 85:20:@8463.4]
  assign _GEN_222 = _T_10325 ? _T_1061_62 : _T_10211_62; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9297.4]
  assign _GEN_223 = _T_10325 ? _T_9253 : _T_10211_63; // @[NV_NVDLA_CSC_WL_dec.scala 104:9:@9302.4]
  assign _T_10413 = _T_10211_0 ? _T_9260_0 : 8'h0; // @[Mux.scala 46:16:@9307.4]
  assign _T_10417 = 2'h2 == _T_10211_1; // @[Mux.scala 46:19:@9309.4]
  assign _T_10418 = _T_10417 ? _T_9260_1 : 8'h0; // @[Mux.scala 46:16:@9310.4]
  assign _T_10419 = 2'h1 == _T_10211_1; // @[Mux.scala 46:19:@9311.4]
  assign _T_10420 = _T_10419 ? _T_9260_0 : _T_10418; // @[Mux.scala 46:16:@9312.4]
  assign _T_10425 = 2'h3 == _T_10211_2; // @[Mux.scala 46:19:@9314.4]
  assign _T_10426 = _T_10425 ? _T_9260_2 : 8'h0; // @[Mux.scala 46:16:@9315.4]
  assign _T_10427 = 2'h2 == _T_10211_2; // @[Mux.scala 46:19:@9316.4]
  assign _T_10428 = _T_10427 ? _T_9260_1 : _T_10426; // @[Mux.scala 46:16:@9317.4]
  assign _T_10429 = 2'h1 == _T_10211_2; // @[Mux.scala 46:19:@9318.4]
  assign _T_10430 = _T_10429 ? _T_9260_0 : _T_10428; // @[Mux.scala 46:16:@9319.4]
  assign _T_10436 = 3'h4 == _T_10211_3; // @[Mux.scala 46:19:@9321.4]
  assign _T_10437 = _T_10436 ? _T_9260_3 : 8'h0; // @[Mux.scala 46:16:@9322.4]
  assign _T_10438 = 3'h3 == _T_10211_3; // @[Mux.scala 46:19:@9323.4]
  assign _T_10439 = _T_10438 ? _T_9260_2 : _T_10437; // @[Mux.scala 46:16:@9324.4]
  assign _T_10440 = 3'h2 == _T_10211_3; // @[Mux.scala 46:19:@9325.4]
  assign _T_10441 = _T_10440 ? _T_9260_1 : _T_10439; // @[Mux.scala 46:16:@9326.4]
  assign _T_10442 = 3'h1 == _T_10211_3; // @[Mux.scala 46:19:@9327.4]
  assign _T_10443 = _T_10442 ? _T_9260_0 : _T_10441; // @[Mux.scala 46:16:@9328.4]
  assign _T_10450 = 3'h5 == _T_10211_4; // @[Mux.scala 46:19:@9330.4]
  assign _T_10451 = _T_10450 ? _T_9260_4 : 8'h0; // @[Mux.scala 46:16:@9331.4]
  assign _T_10452 = 3'h4 == _T_10211_4; // @[Mux.scala 46:19:@9332.4]
  assign _T_10453 = _T_10452 ? _T_9260_3 : _T_10451; // @[Mux.scala 46:16:@9333.4]
  assign _T_10454 = 3'h3 == _T_10211_4; // @[Mux.scala 46:19:@9334.4]
  assign _T_10455 = _T_10454 ? _T_9260_2 : _T_10453; // @[Mux.scala 46:16:@9335.4]
  assign _T_10456 = 3'h2 == _T_10211_4; // @[Mux.scala 46:19:@9336.4]
  assign _T_10457 = _T_10456 ? _T_9260_1 : _T_10455; // @[Mux.scala 46:16:@9337.4]
  assign _T_10458 = 3'h1 == _T_10211_4; // @[Mux.scala 46:19:@9338.4]
  assign _T_10459 = _T_10458 ? _T_9260_0 : _T_10457; // @[Mux.scala 46:16:@9339.4]
  assign _T_10467 = 3'h6 == _T_10211_5; // @[Mux.scala 46:19:@9341.4]
  assign _T_10468 = _T_10467 ? _T_9260_5 : 8'h0; // @[Mux.scala 46:16:@9342.4]
  assign _T_10469 = 3'h5 == _T_10211_5; // @[Mux.scala 46:19:@9343.4]
  assign _T_10470 = _T_10469 ? _T_9260_4 : _T_10468; // @[Mux.scala 46:16:@9344.4]
  assign _T_10471 = 3'h4 == _T_10211_5; // @[Mux.scala 46:19:@9345.4]
  assign _T_10472 = _T_10471 ? _T_9260_3 : _T_10470; // @[Mux.scala 46:16:@9346.4]
  assign _T_10473 = 3'h3 == _T_10211_5; // @[Mux.scala 46:19:@9347.4]
  assign _T_10474 = _T_10473 ? _T_9260_2 : _T_10472; // @[Mux.scala 46:16:@9348.4]
  assign _T_10475 = 3'h2 == _T_10211_5; // @[Mux.scala 46:19:@9349.4]
  assign _T_10476 = _T_10475 ? _T_9260_1 : _T_10474; // @[Mux.scala 46:16:@9350.4]
  assign _T_10477 = 3'h1 == _T_10211_5; // @[Mux.scala 46:19:@9351.4]
  assign _T_10478 = _T_10477 ? _T_9260_0 : _T_10476; // @[Mux.scala 46:16:@9352.4]
  assign _T_10487 = 3'h7 == _T_10211_6; // @[Mux.scala 46:19:@9354.4]
  assign _T_10488 = _T_10487 ? _T_9260_6 : 8'h0; // @[Mux.scala 46:16:@9355.4]
  assign _T_10489 = 3'h6 == _T_10211_6; // @[Mux.scala 46:19:@9356.4]
  assign _T_10490 = _T_10489 ? _T_9260_5 : _T_10488; // @[Mux.scala 46:16:@9357.4]
  assign _T_10491 = 3'h5 == _T_10211_6; // @[Mux.scala 46:19:@9358.4]
  assign _T_10492 = _T_10491 ? _T_9260_4 : _T_10490; // @[Mux.scala 46:16:@9359.4]
  assign _T_10493 = 3'h4 == _T_10211_6; // @[Mux.scala 46:19:@9360.4]
  assign _T_10494 = _T_10493 ? _T_9260_3 : _T_10492; // @[Mux.scala 46:16:@9361.4]
  assign _T_10495 = 3'h3 == _T_10211_6; // @[Mux.scala 46:19:@9362.4]
  assign _T_10496 = _T_10495 ? _T_9260_2 : _T_10494; // @[Mux.scala 46:16:@9363.4]
  assign _T_10497 = 3'h2 == _T_10211_6; // @[Mux.scala 46:19:@9364.4]
  assign _T_10498 = _T_10497 ? _T_9260_1 : _T_10496; // @[Mux.scala 46:16:@9365.4]
  assign _T_10499 = 3'h1 == _T_10211_6; // @[Mux.scala 46:19:@9366.4]
  assign _T_10500 = _T_10499 ? _T_9260_0 : _T_10498; // @[Mux.scala 46:16:@9367.4]
  assign _T_10510 = 4'h8 == _T_10211_7; // @[Mux.scala 46:19:@9369.4]
  assign _T_10511 = _T_10510 ? _T_9260_7 : 8'h0; // @[Mux.scala 46:16:@9370.4]
  assign _T_10512 = 4'h7 == _T_10211_7; // @[Mux.scala 46:19:@9371.4]
  assign _T_10513 = _T_10512 ? _T_9260_6 : _T_10511; // @[Mux.scala 46:16:@9372.4]
  assign _T_10514 = 4'h6 == _T_10211_7; // @[Mux.scala 46:19:@9373.4]
  assign _T_10515 = _T_10514 ? _T_9260_5 : _T_10513; // @[Mux.scala 46:16:@9374.4]
  assign _T_10516 = 4'h5 == _T_10211_7; // @[Mux.scala 46:19:@9375.4]
  assign _T_10517 = _T_10516 ? _T_9260_4 : _T_10515; // @[Mux.scala 46:16:@9376.4]
  assign _T_10518 = 4'h4 == _T_10211_7; // @[Mux.scala 46:19:@9377.4]
  assign _T_10519 = _T_10518 ? _T_9260_3 : _T_10517; // @[Mux.scala 46:16:@9378.4]
  assign _T_10520 = 4'h3 == _T_10211_7; // @[Mux.scala 46:19:@9379.4]
  assign _T_10521 = _T_10520 ? _T_9260_2 : _T_10519; // @[Mux.scala 46:16:@9380.4]
  assign _T_10522 = 4'h2 == _T_10211_7; // @[Mux.scala 46:19:@9381.4]
  assign _T_10523 = _T_10522 ? _T_9260_1 : _T_10521; // @[Mux.scala 46:16:@9382.4]
  assign _T_10524 = 4'h1 == _T_10211_7; // @[Mux.scala 46:19:@9383.4]
  assign _T_10525 = _T_10524 ? _T_9260_0 : _T_10523; // @[Mux.scala 46:16:@9384.4]
  assign _T_10536 = 4'h9 == _T_10211_8; // @[Mux.scala 46:19:@9386.4]
  assign _T_10537 = _T_10536 ? _T_9260_8 : 8'h0; // @[Mux.scala 46:16:@9387.4]
  assign _T_10538 = 4'h8 == _T_10211_8; // @[Mux.scala 46:19:@9388.4]
  assign _T_10539 = _T_10538 ? _T_9260_7 : _T_10537; // @[Mux.scala 46:16:@9389.4]
  assign _T_10540 = 4'h7 == _T_10211_8; // @[Mux.scala 46:19:@9390.4]
  assign _T_10541 = _T_10540 ? _T_9260_6 : _T_10539; // @[Mux.scala 46:16:@9391.4]
  assign _T_10542 = 4'h6 == _T_10211_8; // @[Mux.scala 46:19:@9392.4]
  assign _T_10543 = _T_10542 ? _T_9260_5 : _T_10541; // @[Mux.scala 46:16:@9393.4]
  assign _T_10544 = 4'h5 == _T_10211_8; // @[Mux.scala 46:19:@9394.4]
  assign _T_10545 = _T_10544 ? _T_9260_4 : _T_10543; // @[Mux.scala 46:16:@9395.4]
  assign _T_10546 = 4'h4 == _T_10211_8; // @[Mux.scala 46:19:@9396.4]
  assign _T_10547 = _T_10546 ? _T_9260_3 : _T_10545; // @[Mux.scala 46:16:@9397.4]
  assign _T_10548 = 4'h3 == _T_10211_8; // @[Mux.scala 46:19:@9398.4]
  assign _T_10549 = _T_10548 ? _T_9260_2 : _T_10547; // @[Mux.scala 46:16:@9399.4]
  assign _T_10550 = 4'h2 == _T_10211_8; // @[Mux.scala 46:19:@9400.4]
  assign _T_10551 = _T_10550 ? _T_9260_1 : _T_10549; // @[Mux.scala 46:16:@9401.4]
  assign _T_10552 = 4'h1 == _T_10211_8; // @[Mux.scala 46:19:@9402.4]
  assign _T_10553 = _T_10552 ? _T_9260_0 : _T_10551; // @[Mux.scala 46:16:@9403.4]
  assign _T_10565 = 4'ha == _T_10211_9; // @[Mux.scala 46:19:@9405.4]
  assign _T_10566 = _T_10565 ? _T_9260_9 : 8'h0; // @[Mux.scala 46:16:@9406.4]
  assign _T_10567 = 4'h9 == _T_10211_9; // @[Mux.scala 46:19:@9407.4]
  assign _T_10568 = _T_10567 ? _T_9260_8 : _T_10566; // @[Mux.scala 46:16:@9408.4]
  assign _T_10569 = 4'h8 == _T_10211_9; // @[Mux.scala 46:19:@9409.4]
  assign _T_10570 = _T_10569 ? _T_9260_7 : _T_10568; // @[Mux.scala 46:16:@9410.4]
  assign _T_10571 = 4'h7 == _T_10211_9; // @[Mux.scala 46:19:@9411.4]
  assign _T_10572 = _T_10571 ? _T_9260_6 : _T_10570; // @[Mux.scala 46:16:@9412.4]
  assign _T_10573 = 4'h6 == _T_10211_9; // @[Mux.scala 46:19:@9413.4]
  assign _T_10574 = _T_10573 ? _T_9260_5 : _T_10572; // @[Mux.scala 46:16:@9414.4]
  assign _T_10575 = 4'h5 == _T_10211_9; // @[Mux.scala 46:19:@9415.4]
  assign _T_10576 = _T_10575 ? _T_9260_4 : _T_10574; // @[Mux.scala 46:16:@9416.4]
  assign _T_10577 = 4'h4 == _T_10211_9; // @[Mux.scala 46:19:@9417.4]
  assign _T_10578 = _T_10577 ? _T_9260_3 : _T_10576; // @[Mux.scala 46:16:@9418.4]
  assign _T_10579 = 4'h3 == _T_10211_9; // @[Mux.scala 46:19:@9419.4]
  assign _T_10580 = _T_10579 ? _T_9260_2 : _T_10578; // @[Mux.scala 46:16:@9420.4]
  assign _T_10581 = 4'h2 == _T_10211_9; // @[Mux.scala 46:19:@9421.4]
  assign _T_10582 = _T_10581 ? _T_9260_1 : _T_10580; // @[Mux.scala 46:16:@9422.4]
  assign _T_10583 = 4'h1 == _T_10211_9; // @[Mux.scala 46:19:@9423.4]
  assign _T_10584 = _T_10583 ? _T_9260_0 : _T_10582; // @[Mux.scala 46:16:@9424.4]
  assign _T_10597 = 4'hb == _T_10211_10; // @[Mux.scala 46:19:@9426.4]
  assign _T_10598 = _T_10597 ? _T_9260_10 : 8'h0; // @[Mux.scala 46:16:@9427.4]
  assign _T_10599 = 4'ha == _T_10211_10; // @[Mux.scala 46:19:@9428.4]
  assign _T_10600 = _T_10599 ? _T_9260_9 : _T_10598; // @[Mux.scala 46:16:@9429.4]
  assign _T_10601 = 4'h9 == _T_10211_10; // @[Mux.scala 46:19:@9430.4]
  assign _T_10602 = _T_10601 ? _T_9260_8 : _T_10600; // @[Mux.scala 46:16:@9431.4]
  assign _T_10603 = 4'h8 == _T_10211_10; // @[Mux.scala 46:19:@9432.4]
  assign _T_10604 = _T_10603 ? _T_9260_7 : _T_10602; // @[Mux.scala 46:16:@9433.4]
  assign _T_10605 = 4'h7 == _T_10211_10; // @[Mux.scala 46:19:@9434.4]
  assign _T_10606 = _T_10605 ? _T_9260_6 : _T_10604; // @[Mux.scala 46:16:@9435.4]
  assign _T_10607 = 4'h6 == _T_10211_10; // @[Mux.scala 46:19:@9436.4]
  assign _T_10608 = _T_10607 ? _T_9260_5 : _T_10606; // @[Mux.scala 46:16:@9437.4]
  assign _T_10609 = 4'h5 == _T_10211_10; // @[Mux.scala 46:19:@9438.4]
  assign _T_10610 = _T_10609 ? _T_9260_4 : _T_10608; // @[Mux.scala 46:16:@9439.4]
  assign _T_10611 = 4'h4 == _T_10211_10; // @[Mux.scala 46:19:@9440.4]
  assign _T_10612 = _T_10611 ? _T_9260_3 : _T_10610; // @[Mux.scala 46:16:@9441.4]
  assign _T_10613 = 4'h3 == _T_10211_10; // @[Mux.scala 46:19:@9442.4]
  assign _T_10614 = _T_10613 ? _T_9260_2 : _T_10612; // @[Mux.scala 46:16:@9443.4]
  assign _T_10615 = 4'h2 == _T_10211_10; // @[Mux.scala 46:19:@9444.4]
  assign _T_10616 = _T_10615 ? _T_9260_1 : _T_10614; // @[Mux.scala 46:16:@9445.4]
  assign _T_10617 = 4'h1 == _T_10211_10; // @[Mux.scala 46:19:@9446.4]
  assign _T_10618 = _T_10617 ? _T_9260_0 : _T_10616; // @[Mux.scala 46:16:@9447.4]
  assign _T_10632 = 4'hc == _T_10211_11; // @[Mux.scala 46:19:@9449.4]
  assign _T_10633 = _T_10632 ? _T_9260_11 : 8'h0; // @[Mux.scala 46:16:@9450.4]
  assign _T_10634 = 4'hb == _T_10211_11; // @[Mux.scala 46:19:@9451.4]
  assign _T_10635 = _T_10634 ? _T_9260_10 : _T_10633; // @[Mux.scala 46:16:@9452.4]
  assign _T_10636 = 4'ha == _T_10211_11; // @[Mux.scala 46:19:@9453.4]
  assign _T_10637 = _T_10636 ? _T_9260_9 : _T_10635; // @[Mux.scala 46:16:@9454.4]
  assign _T_10638 = 4'h9 == _T_10211_11; // @[Mux.scala 46:19:@9455.4]
  assign _T_10639 = _T_10638 ? _T_9260_8 : _T_10637; // @[Mux.scala 46:16:@9456.4]
  assign _T_10640 = 4'h8 == _T_10211_11; // @[Mux.scala 46:19:@9457.4]
  assign _T_10641 = _T_10640 ? _T_9260_7 : _T_10639; // @[Mux.scala 46:16:@9458.4]
  assign _T_10642 = 4'h7 == _T_10211_11; // @[Mux.scala 46:19:@9459.4]
  assign _T_10643 = _T_10642 ? _T_9260_6 : _T_10641; // @[Mux.scala 46:16:@9460.4]
  assign _T_10644 = 4'h6 == _T_10211_11; // @[Mux.scala 46:19:@9461.4]
  assign _T_10645 = _T_10644 ? _T_9260_5 : _T_10643; // @[Mux.scala 46:16:@9462.4]
  assign _T_10646 = 4'h5 == _T_10211_11; // @[Mux.scala 46:19:@9463.4]
  assign _T_10647 = _T_10646 ? _T_9260_4 : _T_10645; // @[Mux.scala 46:16:@9464.4]
  assign _T_10648 = 4'h4 == _T_10211_11; // @[Mux.scala 46:19:@9465.4]
  assign _T_10649 = _T_10648 ? _T_9260_3 : _T_10647; // @[Mux.scala 46:16:@9466.4]
  assign _T_10650 = 4'h3 == _T_10211_11; // @[Mux.scala 46:19:@9467.4]
  assign _T_10651 = _T_10650 ? _T_9260_2 : _T_10649; // @[Mux.scala 46:16:@9468.4]
  assign _T_10652 = 4'h2 == _T_10211_11; // @[Mux.scala 46:19:@9469.4]
  assign _T_10653 = _T_10652 ? _T_9260_1 : _T_10651; // @[Mux.scala 46:16:@9470.4]
  assign _T_10654 = 4'h1 == _T_10211_11; // @[Mux.scala 46:19:@9471.4]
  assign _T_10655 = _T_10654 ? _T_9260_0 : _T_10653; // @[Mux.scala 46:16:@9472.4]
  assign _T_10670 = 4'hd == _T_10211_12; // @[Mux.scala 46:19:@9474.4]
  assign _T_10671 = _T_10670 ? _T_9260_12 : 8'h0; // @[Mux.scala 46:16:@9475.4]
  assign _T_10672 = 4'hc == _T_10211_12; // @[Mux.scala 46:19:@9476.4]
  assign _T_10673 = _T_10672 ? _T_9260_11 : _T_10671; // @[Mux.scala 46:16:@9477.4]
  assign _T_10674 = 4'hb == _T_10211_12; // @[Mux.scala 46:19:@9478.4]
  assign _T_10675 = _T_10674 ? _T_9260_10 : _T_10673; // @[Mux.scala 46:16:@9479.4]
  assign _T_10676 = 4'ha == _T_10211_12; // @[Mux.scala 46:19:@9480.4]
  assign _T_10677 = _T_10676 ? _T_9260_9 : _T_10675; // @[Mux.scala 46:16:@9481.4]
  assign _T_10678 = 4'h9 == _T_10211_12; // @[Mux.scala 46:19:@9482.4]
  assign _T_10679 = _T_10678 ? _T_9260_8 : _T_10677; // @[Mux.scala 46:16:@9483.4]
  assign _T_10680 = 4'h8 == _T_10211_12; // @[Mux.scala 46:19:@9484.4]
  assign _T_10681 = _T_10680 ? _T_9260_7 : _T_10679; // @[Mux.scala 46:16:@9485.4]
  assign _T_10682 = 4'h7 == _T_10211_12; // @[Mux.scala 46:19:@9486.4]
  assign _T_10683 = _T_10682 ? _T_9260_6 : _T_10681; // @[Mux.scala 46:16:@9487.4]
  assign _T_10684 = 4'h6 == _T_10211_12; // @[Mux.scala 46:19:@9488.4]
  assign _T_10685 = _T_10684 ? _T_9260_5 : _T_10683; // @[Mux.scala 46:16:@9489.4]
  assign _T_10686 = 4'h5 == _T_10211_12; // @[Mux.scala 46:19:@9490.4]
  assign _T_10687 = _T_10686 ? _T_9260_4 : _T_10685; // @[Mux.scala 46:16:@9491.4]
  assign _T_10688 = 4'h4 == _T_10211_12; // @[Mux.scala 46:19:@9492.4]
  assign _T_10689 = _T_10688 ? _T_9260_3 : _T_10687; // @[Mux.scala 46:16:@9493.4]
  assign _T_10690 = 4'h3 == _T_10211_12; // @[Mux.scala 46:19:@9494.4]
  assign _T_10691 = _T_10690 ? _T_9260_2 : _T_10689; // @[Mux.scala 46:16:@9495.4]
  assign _T_10692 = 4'h2 == _T_10211_12; // @[Mux.scala 46:19:@9496.4]
  assign _T_10693 = _T_10692 ? _T_9260_1 : _T_10691; // @[Mux.scala 46:16:@9497.4]
  assign _T_10694 = 4'h1 == _T_10211_12; // @[Mux.scala 46:19:@9498.4]
  assign _T_10695 = _T_10694 ? _T_9260_0 : _T_10693; // @[Mux.scala 46:16:@9499.4]
  assign _T_10711 = 4'he == _T_10211_13; // @[Mux.scala 46:19:@9501.4]
  assign _T_10712 = _T_10711 ? _T_9260_13 : 8'h0; // @[Mux.scala 46:16:@9502.4]
  assign _T_10713 = 4'hd == _T_10211_13; // @[Mux.scala 46:19:@9503.4]
  assign _T_10714 = _T_10713 ? _T_9260_12 : _T_10712; // @[Mux.scala 46:16:@9504.4]
  assign _T_10715 = 4'hc == _T_10211_13; // @[Mux.scala 46:19:@9505.4]
  assign _T_10716 = _T_10715 ? _T_9260_11 : _T_10714; // @[Mux.scala 46:16:@9506.4]
  assign _T_10717 = 4'hb == _T_10211_13; // @[Mux.scala 46:19:@9507.4]
  assign _T_10718 = _T_10717 ? _T_9260_10 : _T_10716; // @[Mux.scala 46:16:@9508.4]
  assign _T_10719 = 4'ha == _T_10211_13; // @[Mux.scala 46:19:@9509.4]
  assign _T_10720 = _T_10719 ? _T_9260_9 : _T_10718; // @[Mux.scala 46:16:@9510.4]
  assign _T_10721 = 4'h9 == _T_10211_13; // @[Mux.scala 46:19:@9511.4]
  assign _T_10722 = _T_10721 ? _T_9260_8 : _T_10720; // @[Mux.scala 46:16:@9512.4]
  assign _T_10723 = 4'h8 == _T_10211_13; // @[Mux.scala 46:19:@9513.4]
  assign _T_10724 = _T_10723 ? _T_9260_7 : _T_10722; // @[Mux.scala 46:16:@9514.4]
  assign _T_10725 = 4'h7 == _T_10211_13; // @[Mux.scala 46:19:@9515.4]
  assign _T_10726 = _T_10725 ? _T_9260_6 : _T_10724; // @[Mux.scala 46:16:@9516.4]
  assign _T_10727 = 4'h6 == _T_10211_13; // @[Mux.scala 46:19:@9517.4]
  assign _T_10728 = _T_10727 ? _T_9260_5 : _T_10726; // @[Mux.scala 46:16:@9518.4]
  assign _T_10729 = 4'h5 == _T_10211_13; // @[Mux.scala 46:19:@9519.4]
  assign _T_10730 = _T_10729 ? _T_9260_4 : _T_10728; // @[Mux.scala 46:16:@9520.4]
  assign _T_10731 = 4'h4 == _T_10211_13; // @[Mux.scala 46:19:@9521.4]
  assign _T_10732 = _T_10731 ? _T_9260_3 : _T_10730; // @[Mux.scala 46:16:@9522.4]
  assign _T_10733 = 4'h3 == _T_10211_13; // @[Mux.scala 46:19:@9523.4]
  assign _T_10734 = _T_10733 ? _T_9260_2 : _T_10732; // @[Mux.scala 46:16:@9524.4]
  assign _T_10735 = 4'h2 == _T_10211_13; // @[Mux.scala 46:19:@9525.4]
  assign _T_10736 = _T_10735 ? _T_9260_1 : _T_10734; // @[Mux.scala 46:16:@9526.4]
  assign _T_10737 = 4'h1 == _T_10211_13; // @[Mux.scala 46:19:@9527.4]
  assign _T_10738 = _T_10737 ? _T_9260_0 : _T_10736; // @[Mux.scala 46:16:@9528.4]
  assign _T_10755 = 4'hf == _T_10211_14; // @[Mux.scala 46:19:@9530.4]
  assign _T_10756 = _T_10755 ? _T_9260_14 : 8'h0; // @[Mux.scala 46:16:@9531.4]
  assign _T_10757 = 4'he == _T_10211_14; // @[Mux.scala 46:19:@9532.4]
  assign _T_10758 = _T_10757 ? _T_9260_13 : _T_10756; // @[Mux.scala 46:16:@9533.4]
  assign _T_10759 = 4'hd == _T_10211_14; // @[Mux.scala 46:19:@9534.4]
  assign _T_10760 = _T_10759 ? _T_9260_12 : _T_10758; // @[Mux.scala 46:16:@9535.4]
  assign _T_10761 = 4'hc == _T_10211_14; // @[Mux.scala 46:19:@9536.4]
  assign _T_10762 = _T_10761 ? _T_9260_11 : _T_10760; // @[Mux.scala 46:16:@9537.4]
  assign _T_10763 = 4'hb == _T_10211_14; // @[Mux.scala 46:19:@9538.4]
  assign _T_10764 = _T_10763 ? _T_9260_10 : _T_10762; // @[Mux.scala 46:16:@9539.4]
  assign _T_10765 = 4'ha == _T_10211_14; // @[Mux.scala 46:19:@9540.4]
  assign _T_10766 = _T_10765 ? _T_9260_9 : _T_10764; // @[Mux.scala 46:16:@9541.4]
  assign _T_10767 = 4'h9 == _T_10211_14; // @[Mux.scala 46:19:@9542.4]
  assign _T_10768 = _T_10767 ? _T_9260_8 : _T_10766; // @[Mux.scala 46:16:@9543.4]
  assign _T_10769 = 4'h8 == _T_10211_14; // @[Mux.scala 46:19:@9544.4]
  assign _T_10770 = _T_10769 ? _T_9260_7 : _T_10768; // @[Mux.scala 46:16:@9545.4]
  assign _T_10771 = 4'h7 == _T_10211_14; // @[Mux.scala 46:19:@9546.4]
  assign _T_10772 = _T_10771 ? _T_9260_6 : _T_10770; // @[Mux.scala 46:16:@9547.4]
  assign _T_10773 = 4'h6 == _T_10211_14; // @[Mux.scala 46:19:@9548.4]
  assign _T_10774 = _T_10773 ? _T_9260_5 : _T_10772; // @[Mux.scala 46:16:@9549.4]
  assign _T_10775 = 4'h5 == _T_10211_14; // @[Mux.scala 46:19:@9550.4]
  assign _T_10776 = _T_10775 ? _T_9260_4 : _T_10774; // @[Mux.scala 46:16:@9551.4]
  assign _T_10777 = 4'h4 == _T_10211_14; // @[Mux.scala 46:19:@9552.4]
  assign _T_10778 = _T_10777 ? _T_9260_3 : _T_10776; // @[Mux.scala 46:16:@9553.4]
  assign _T_10779 = 4'h3 == _T_10211_14; // @[Mux.scala 46:19:@9554.4]
  assign _T_10780 = _T_10779 ? _T_9260_2 : _T_10778; // @[Mux.scala 46:16:@9555.4]
  assign _T_10781 = 4'h2 == _T_10211_14; // @[Mux.scala 46:19:@9556.4]
  assign _T_10782 = _T_10781 ? _T_9260_1 : _T_10780; // @[Mux.scala 46:16:@9557.4]
  assign _T_10783 = 4'h1 == _T_10211_14; // @[Mux.scala 46:19:@9558.4]
  assign _T_10784 = _T_10783 ? _T_9260_0 : _T_10782; // @[Mux.scala 46:16:@9559.4]
  assign _T_10802 = 5'h10 == _T_10211_15; // @[Mux.scala 46:19:@9561.4]
  assign _T_10803 = _T_10802 ? _T_9260_15 : 8'h0; // @[Mux.scala 46:16:@9562.4]
  assign _T_10804 = 5'hf == _T_10211_15; // @[Mux.scala 46:19:@9563.4]
  assign _T_10805 = _T_10804 ? _T_9260_14 : _T_10803; // @[Mux.scala 46:16:@9564.4]
  assign _T_10806 = 5'he == _T_10211_15; // @[Mux.scala 46:19:@9565.4]
  assign _T_10807 = _T_10806 ? _T_9260_13 : _T_10805; // @[Mux.scala 46:16:@9566.4]
  assign _T_10808 = 5'hd == _T_10211_15; // @[Mux.scala 46:19:@9567.4]
  assign _T_10809 = _T_10808 ? _T_9260_12 : _T_10807; // @[Mux.scala 46:16:@9568.4]
  assign _T_10810 = 5'hc == _T_10211_15; // @[Mux.scala 46:19:@9569.4]
  assign _T_10811 = _T_10810 ? _T_9260_11 : _T_10809; // @[Mux.scala 46:16:@9570.4]
  assign _T_10812 = 5'hb == _T_10211_15; // @[Mux.scala 46:19:@9571.4]
  assign _T_10813 = _T_10812 ? _T_9260_10 : _T_10811; // @[Mux.scala 46:16:@9572.4]
  assign _T_10814 = 5'ha == _T_10211_15; // @[Mux.scala 46:19:@9573.4]
  assign _T_10815 = _T_10814 ? _T_9260_9 : _T_10813; // @[Mux.scala 46:16:@9574.4]
  assign _T_10816 = 5'h9 == _T_10211_15; // @[Mux.scala 46:19:@9575.4]
  assign _T_10817 = _T_10816 ? _T_9260_8 : _T_10815; // @[Mux.scala 46:16:@9576.4]
  assign _T_10818 = 5'h8 == _T_10211_15; // @[Mux.scala 46:19:@9577.4]
  assign _T_10819 = _T_10818 ? _T_9260_7 : _T_10817; // @[Mux.scala 46:16:@9578.4]
  assign _T_10820 = 5'h7 == _T_10211_15; // @[Mux.scala 46:19:@9579.4]
  assign _T_10821 = _T_10820 ? _T_9260_6 : _T_10819; // @[Mux.scala 46:16:@9580.4]
  assign _T_10822 = 5'h6 == _T_10211_15; // @[Mux.scala 46:19:@9581.4]
  assign _T_10823 = _T_10822 ? _T_9260_5 : _T_10821; // @[Mux.scala 46:16:@9582.4]
  assign _T_10824 = 5'h5 == _T_10211_15; // @[Mux.scala 46:19:@9583.4]
  assign _T_10825 = _T_10824 ? _T_9260_4 : _T_10823; // @[Mux.scala 46:16:@9584.4]
  assign _T_10826 = 5'h4 == _T_10211_15; // @[Mux.scala 46:19:@9585.4]
  assign _T_10827 = _T_10826 ? _T_9260_3 : _T_10825; // @[Mux.scala 46:16:@9586.4]
  assign _T_10828 = 5'h3 == _T_10211_15; // @[Mux.scala 46:19:@9587.4]
  assign _T_10829 = _T_10828 ? _T_9260_2 : _T_10827; // @[Mux.scala 46:16:@9588.4]
  assign _T_10830 = 5'h2 == _T_10211_15; // @[Mux.scala 46:19:@9589.4]
  assign _T_10831 = _T_10830 ? _T_9260_1 : _T_10829; // @[Mux.scala 46:16:@9590.4]
  assign _T_10832 = 5'h1 == _T_10211_15; // @[Mux.scala 46:19:@9591.4]
  assign _T_10833 = _T_10832 ? _T_9260_0 : _T_10831; // @[Mux.scala 46:16:@9592.4]
  assign _T_10852 = 5'h11 == _T_10211_16; // @[Mux.scala 46:19:@9594.4]
  assign _T_10853 = _T_10852 ? _T_9260_16 : 8'h0; // @[Mux.scala 46:16:@9595.4]
  assign _T_10854 = 5'h10 == _T_10211_16; // @[Mux.scala 46:19:@9596.4]
  assign _T_10855 = _T_10854 ? _T_9260_15 : _T_10853; // @[Mux.scala 46:16:@9597.4]
  assign _T_10856 = 5'hf == _T_10211_16; // @[Mux.scala 46:19:@9598.4]
  assign _T_10857 = _T_10856 ? _T_9260_14 : _T_10855; // @[Mux.scala 46:16:@9599.4]
  assign _T_10858 = 5'he == _T_10211_16; // @[Mux.scala 46:19:@9600.4]
  assign _T_10859 = _T_10858 ? _T_9260_13 : _T_10857; // @[Mux.scala 46:16:@9601.4]
  assign _T_10860 = 5'hd == _T_10211_16; // @[Mux.scala 46:19:@9602.4]
  assign _T_10861 = _T_10860 ? _T_9260_12 : _T_10859; // @[Mux.scala 46:16:@9603.4]
  assign _T_10862 = 5'hc == _T_10211_16; // @[Mux.scala 46:19:@9604.4]
  assign _T_10863 = _T_10862 ? _T_9260_11 : _T_10861; // @[Mux.scala 46:16:@9605.4]
  assign _T_10864 = 5'hb == _T_10211_16; // @[Mux.scala 46:19:@9606.4]
  assign _T_10865 = _T_10864 ? _T_9260_10 : _T_10863; // @[Mux.scala 46:16:@9607.4]
  assign _T_10866 = 5'ha == _T_10211_16; // @[Mux.scala 46:19:@9608.4]
  assign _T_10867 = _T_10866 ? _T_9260_9 : _T_10865; // @[Mux.scala 46:16:@9609.4]
  assign _T_10868 = 5'h9 == _T_10211_16; // @[Mux.scala 46:19:@9610.4]
  assign _T_10869 = _T_10868 ? _T_9260_8 : _T_10867; // @[Mux.scala 46:16:@9611.4]
  assign _T_10870 = 5'h8 == _T_10211_16; // @[Mux.scala 46:19:@9612.4]
  assign _T_10871 = _T_10870 ? _T_9260_7 : _T_10869; // @[Mux.scala 46:16:@9613.4]
  assign _T_10872 = 5'h7 == _T_10211_16; // @[Mux.scala 46:19:@9614.4]
  assign _T_10873 = _T_10872 ? _T_9260_6 : _T_10871; // @[Mux.scala 46:16:@9615.4]
  assign _T_10874 = 5'h6 == _T_10211_16; // @[Mux.scala 46:19:@9616.4]
  assign _T_10875 = _T_10874 ? _T_9260_5 : _T_10873; // @[Mux.scala 46:16:@9617.4]
  assign _T_10876 = 5'h5 == _T_10211_16; // @[Mux.scala 46:19:@9618.4]
  assign _T_10877 = _T_10876 ? _T_9260_4 : _T_10875; // @[Mux.scala 46:16:@9619.4]
  assign _T_10878 = 5'h4 == _T_10211_16; // @[Mux.scala 46:19:@9620.4]
  assign _T_10879 = _T_10878 ? _T_9260_3 : _T_10877; // @[Mux.scala 46:16:@9621.4]
  assign _T_10880 = 5'h3 == _T_10211_16; // @[Mux.scala 46:19:@9622.4]
  assign _T_10881 = _T_10880 ? _T_9260_2 : _T_10879; // @[Mux.scala 46:16:@9623.4]
  assign _T_10882 = 5'h2 == _T_10211_16; // @[Mux.scala 46:19:@9624.4]
  assign _T_10883 = _T_10882 ? _T_9260_1 : _T_10881; // @[Mux.scala 46:16:@9625.4]
  assign _T_10884 = 5'h1 == _T_10211_16; // @[Mux.scala 46:19:@9626.4]
  assign _T_10885 = _T_10884 ? _T_9260_0 : _T_10883; // @[Mux.scala 46:16:@9627.4]
  assign _T_10905 = 5'h12 == _T_10211_17; // @[Mux.scala 46:19:@9629.4]
  assign _T_10906 = _T_10905 ? _T_9260_17 : 8'h0; // @[Mux.scala 46:16:@9630.4]
  assign _T_10907 = 5'h11 == _T_10211_17; // @[Mux.scala 46:19:@9631.4]
  assign _T_10908 = _T_10907 ? _T_9260_16 : _T_10906; // @[Mux.scala 46:16:@9632.4]
  assign _T_10909 = 5'h10 == _T_10211_17; // @[Mux.scala 46:19:@9633.4]
  assign _T_10910 = _T_10909 ? _T_9260_15 : _T_10908; // @[Mux.scala 46:16:@9634.4]
  assign _T_10911 = 5'hf == _T_10211_17; // @[Mux.scala 46:19:@9635.4]
  assign _T_10912 = _T_10911 ? _T_9260_14 : _T_10910; // @[Mux.scala 46:16:@9636.4]
  assign _T_10913 = 5'he == _T_10211_17; // @[Mux.scala 46:19:@9637.4]
  assign _T_10914 = _T_10913 ? _T_9260_13 : _T_10912; // @[Mux.scala 46:16:@9638.4]
  assign _T_10915 = 5'hd == _T_10211_17; // @[Mux.scala 46:19:@9639.4]
  assign _T_10916 = _T_10915 ? _T_9260_12 : _T_10914; // @[Mux.scala 46:16:@9640.4]
  assign _T_10917 = 5'hc == _T_10211_17; // @[Mux.scala 46:19:@9641.4]
  assign _T_10918 = _T_10917 ? _T_9260_11 : _T_10916; // @[Mux.scala 46:16:@9642.4]
  assign _T_10919 = 5'hb == _T_10211_17; // @[Mux.scala 46:19:@9643.4]
  assign _T_10920 = _T_10919 ? _T_9260_10 : _T_10918; // @[Mux.scala 46:16:@9644.4]
  assign _T_10921 = 5'ha == _T_10211_17; // @[Mux.scala 46:19:@9645.4]
  assign _T_10922 = _T_10921 ? _T_9260_9 : _T_10920; // @[Mux.scala 46:16:@9646.4]
  assign _T_10923 = 5'h9 == _T_10211_17; // @[Mux.scala 46:19:@9647.4]
  assign _T_10924 = _T_10923 ? _T_9260_8 : _T_10922; // @[Mux.scala 46:16:@9648.4]
  assign _T_10925 = 5'h8 == _T_10211_17; // @[Mux.scala 46:19:@9649.4]
  assign _T_10926 = _T_10925 ? _T_9260_7 : _T_10924; // @[Mux.scala 46:16:@9650.4]
  assign _T_10927 = 5'h7 == _T_10211_17; // @[Mux.scala 46:19:@9651.4]
  assign _T_10928 = _T_10927 ? _T_9260_6 : _T_10926; // @[Mux.scala 46:16:@9652.4]
  assign _T_10929 = 5'h6 == _T_10211_17; // @[Mux.scala 46:19:@9653.4]
  assign _T_10930 = _T_10929 ? _T_9260_5 : _T_10928; // @[Mux.scala 46:16:@9654.4]
  assign _T_10931 = 5'h5 == _T_10211_17; // @[Mux.scala 46:19:@9655.4]
  assign _T_10932 = _T_10931 ? _T_9260_4 : _T_10930; // @[Mux.scala 46:16:@9656.4]
  assign _T_10933 = 5'h4 == _T_10211_17; // @[Mux.scala 46:19:@9657.4]
  assign _T_10934 = _T_10933 ? _T_9260_3 : _T_10932; // @[Mux.scala 46:16:@9658.4]
  assign _T_10935 = 5'h3 == _T_10211_17; // @[Mux.scala 46:19:@9659.4]
  assign _T_10936 = _T_10935 ? _T_9260_2 : _T_10934; // @[Mux.scala 46:16:@9660.4]
  assign _T_10937 = 5'h2 == _T_10211_17; // @[Mux.scala 46:19:@9661.4]
  assign _T_10938 = _T_10937 ? _T_9260_1 : _T_10936; // @[Mux.scala 46:16:@9662.4]
  assign _T_10939 = 5'h1 == _T_10211_17; // @[Mux.scala 46:19:@9663.4]
  assign _T_10940 = _T_10939 ? _T_9260_0 : _T_10938; // @[Mux.scala 46:16:@9664.4]
  assign _T_10961 = 5'h13 == _T_10211_18; // @[Mux.scala 46:19:@9666.4]
  assign _T_10962 = _T_10961 ? _T_9260_18 : 8'h0; // @[Mux.scala 46:16:@9667.4]
  assign _T_10963 = 5'h12 == _T_10211_18; // @[Mux.scala 46:19:@9668.4]
  assign _T_10964 = _T_10963 ? _T_9260_17 : _T_10962; // @[Mux.scala 46:16:@9669.4]
  assign _T_10965 = 5'h11 == _T_10211_18; // @[Mux.scala 46:19:@9670.4]
  assign _T_10966 = _T_10965 ? _T_9260_16 : _T_10964; // @[Mux.scala 46:16:@9671.4]
  assign _T_10967 = 5'h10 == _T_10211_18; // @[Mux.scala 46:19:@9672.4]
  assign _T_10968 = _T_10967 ? _T_9260_15 : _T_10966; // @[Mux.scala 46:16:@9673.4]
  assign _T_10969 = 5'hf == _T_10211_18; // @[Mux.scala 46:19:@9674.4]
  assign _T_10970 = _T_10969 ? _T_9260_14 : _T_10968; // @[Mux.scala 46:16:@9675.4]
  assign _T_10971 = 5'he == _T_10211_18; // @[Mux.scala 46:19:@9676.4]
  assign _T_10972 = _T_10971 ? _T_9260_13 : _T_10970; // @[Mux.scala 46:16:@9677.4]
  assign _T_10973 = 5'hd == _T_10211_18; // @[Mux.scala 46:19:@9678.4]
  assign _T_10974 = _T_10973 ? _T_9260_12 : _T_10972; // @[Mux.scala 46:16:@9679.4]
  assign _T_10975 = 5'hc == _T_10211_18; // @[Mux.scala 46:19:@9680.4]
  assign _T_10976 = _T_10975 ? _T_9260_11 : _T_10974; // @[Mux.scala 46:16:@9681.4]
  assign _T_10977 = 5'hb == _T_10211_18; // @[Mux.scala 46:19:@9682.4]
  assign _T_10978 = _T_10977 ? _T_9260_10 : _T_10976; // @[Mux.scala 46:16:@9683.4]
  assign _T_10979 = 5'ha == _T_10211_18; // @[Mux.scala 46:19:@9684.4]
  assign _T_10980 = _T_10979 ? _T_9260_9 : _T_10978; // @[Mux.scala 46:16:@9685.4]
  assign _T_10981 = 5'h9 == _T_10211_18; // @[Mux.scala 46:19:@9686.4]
  assign _T_10982 = _T_10981 ? _T_9260_8 : _T_10980; // @[Mux.scala 46:16:@9687.4]
  assign _T_10983 = 5'h8 == _T_10211_18; // @[Mux.scala 46:19:@9688.4]
  assign _T_10984 = _T_10983 ? _T_9260_7 : _T_10982; // @[Mux.scala 46:16:@9689.4]
  assign _T_10985 = 5'h7 == _T_10211_18; // @[Mux.scala 46:19:@9690.4]
  assign _T_10986 = _T_10985 ? _T_9260_6 : _T_10984; // @[Mux.scala 46:16:@9691.4]
  assign _T_10987 = 5'h6 == _T_10211_18; // @[Mux.scala 46:19:@9692.4]
  assign _T_10988 = _T_10987 ? _T_9260_5 : _T_10986; // @[Mux.scala 46:16:@9693.4]
  assign _T_10989 = 5'h5 == _T_10211_18; // @[Mux.scala 46:19:@9694.4]
  assign _T_10990 = _T_10989 ? _T_9260_4 : _T_10988; // @[Mux.scala 46:16:@9695.4]
  assign _T_10991 = 5'h4 == _T_10211_18; // @[Mux.scala 46:19:@9696.4]
  assign _T_10992 = _T_10991 ? _T_9260_3 : _T_10990; // @[Mux.scala 46:16:@9697.4]
  assign _T_10993 = 5'h3 == _T_10211_18; // @[Mux.scala 46:19:@9698.4]
  assign _T_10994 = _T_10993 ? _T_9260_2 : _T_10992; // @[Mux.scala 46:16:@9699.4]
  assign _T_10995 = 5'h2 == _T_10211_18; // @[Mux.scala 46:19:@9700.4]
  assign _T_10996 = _T_10995 ? _T_9260_1 : _T_10994; // @[Mux.scala 46:16:@9701.4]
  assign _T_10997 = 5'h1 == _T_10211_18; // @[Mux.scala 46:19:@9702.4]
  assign _T_10998 = _T_10997 ? _T_9260_0 : _T_10996; // @[Mux.scala 46:16:@9703.4]
  assign _T_11020 = 5'h14 == _T_10211_19; // @[Mux.scala 46:19:@9705.4]
  assign _T_11021 = _T_11020 ? _T_9260_19 : 8'h0; // @[Mux.scala 46:16:@9706.4]
  assign _T_11022 = 5'h13 == _T_10211_19; // @[Mux.scala 46:19:@9707.4]
  assign _T_11023 = _T_11022 ? _T_9260_18 : _T_11021; // @[Mux.scala 46:16:@9708.4]
  assign _T_11024 = 5'h12 == _T_10211_19; // @[Mux.scala 46:19:@9709.4]
  assign _T_11025 = _T_11024 ? _T_9260_17 : _T_11023; // @[Mux.scala 46:16:@9710.4]
  assign _T_11026 = 5'h11 == _T_10211_19; // @[Mux.scala 46:19:@9711.4]
  assign _T_11027 = _T_11026 ? _T_9260_16 : _T_11025; // @[Mux.scala 46:16:@9712.4]
  assign _T_11028 = 5'h10 == _T_10211_19; // @[Mux.scala 46:19:@9713.4]
  assign _T_11029 = _T_11028 ? _T_9260_15 : _T_11027; // @[Mux.scala 46:16:@9714.4]
  assign _T_11030 = 5'hf == _T_10211_19; // @[Mux.scala 46:19:@9715.4]
  assign _T_11031 = _T_11030 ? _T_9260_14 : _T_11029; // @[Mux.scala 46:16:@9716.4]
  assign _T_11032 = 5'he == _T_10211_19; // @[Mux.scala 46:19:@9717.4]
  assign _T_11033 = _T_11032 ? _T_9260_13 : _T_11031; // @[Mux.scala 46:16:@9718.4]
  assign _T_11034 = 5'hd == _T_10211_19; // @[Mux.scala 46:19:@9719.4]
  assign _T_11035 = _T_11034 ? _T_9260_12 : _T_11033; // @[Mux.scala 46:16:@9720.4]
  assign _T_11036 = 5'hc == _T_10211_19; // @[Mux.scala 46:19:@9721.4]
  assign _T_11037 = _T_11036 ? _T_9260_11 : _T_11035; // @[Mux.scala 46:16:@9722.4]
  assign _T_11038 = 5'hb == _T_10211_19; // @[Mux.scala 46:19:@9723.4]
  assign _T_11039 = _T_11038 ? _T_9260_10 : _T_11037; // @[Mux.scala 46:16:@9724.4]
  assign _T_11040 = 5'ha == _T_10211_19; // @[Mux.scala 46:19:@9725.4]
  assign _T_11041 = _T_11040 ? _T_9260_9 : _T_11039; // @[Mux.scala 46:16:@9726.4]
  assign _T_11042 = 5'h9 == _T_10211_19; // @[Mux.scala 46:19:@9727.4]
  assign _T_11043 = _T_11042 ? _T_9260_8 : _T_11041; // @[Mux.scala 46:16:@9728.4]
  assign _T_11044 = 5'h8 == _T_10211_19; // @[Mux.scala 46:19:@9729.4]
  assign _T_11045 = _T_11044 ? _T_9260_7 : _T_11043; // @[Mux.scala 46:16:@9730.4]
  assign _T_11046 = 5'h7 == _T_10211_19; // @[Mux.scala 46:19:@9731.4]
  assign _T_11047 = _T_11046 ? _T_9260_6 : _T_11045; // @[Mux.scala 46:16:@9732.4]
  assign _T_11048 = 5'h6 == _T_10211_19; // @[Mux.scala 46:19:@9733.4]
  assign _T_11049 = _T_11048 ? _T_9260_5 : _T_11047; // @[Mux.scala 46:16:@9734.4]
  assign _T_11050 = 5'h5 == _T_10211_19; // @[Mux.scala 46:19:@9735.4]
  assign _T_11051 = _T_11050 ? _T_9260_4 : _T_11049; // @[Mux.scala 46:16:@9736.4]
  assign _T_11052 = 5'h4 == _T_10211_19; // @[Mux.scala 46:19:@9737.4]
  assign _T_11053 = _T_11052 ? _T_9260_3 : _T_11051; // @[Mux.scala 46:16:@9738.4]
  assign _T_11054 = 5'h3 == _T_10211_19; // @[Mux.scala 46:19:@9739.4]
  assign _T_11055 = _T_11054 ? _T_9260_2 : _T_11053; // @[Mux.scala 46:16:@9740.4]
  assign _T_11056 = 5'h2 == _T_10211_19; // @[Mux.scala 46:19:@9741.4]
  assign _T_11057 = _T_11056 ? _T_9260_1 : _T_11055; // @[Mux.scala 46:16:@9742.4]
  assign _T_11058 = 5'h1 == _T_10211_19; // @[Mux.scala 46:19:@9743.4]
  assign _T_11059 = _T_11058 ? _T_9260_0 : _T_11057; // @[Mux.scala 46:16:@9744.4]
  assign _T_11082 = 5'h15 == _T_10211_20; // @[Mux.scala 46:19:@9746.4]
  assign _T_11083 = _T_11082 ? _T_9260_20 : 8'h0; // @[Mux.scala 46:16:@9747.4]
  assign _T_11084 = 5'h14 == _T_10211_20; // @[Mux.scala 46:19:@9748.4]
  assign _T_11085 = _T_11084 ? _T_9260_19 : _T_11083; // @[Mux.scala 46:16:@9749.4]
  assign _T_11086 = 5'h13 == _T_10211_20; // @[Mux.scala 46:19:@9750.4]
  assign _T_11087 = _T_11086 ? _T_9260_18 : _T_11085; // @[Mux.scala 46:16:@9751.4]
  assign _T_11088 = 5'h12 == _T_10211_20; // @[Mux.scala 46:19:@9752.4]
  assign _T_11089 = _T_11088 ? _T_9260_17 : _T_11087; // @[Mux.scala 46:16:@9753.4]
  assign _T_11090 = 5'h11 == _T_10211_20; // @[Mux.scala 46:19:@9754.4]
  assign _T_11091 = _T_11090 ? _T_9260_16 : _T_11089; // @[Mux.scala 46:16:@9755.4]
  assign _T_11092 = 5'h10 == _T_10211_20; // @[Mux.scala 46:19:@9756.4]
  assign _T_11093 = _T_11092 ? _T_9260_15 : _T_11091; // @[Mux.scala 46:16:@9757.4]
  assign _T_11094 = 5'hf == _T_10211_20; // @[Mux.scala 46:19:@9758.4]
  assign _T_11095 = _T_11094 ? _T_9260_14 : _T_11093; // @[Mux.scala 46:16:@9759.4]
  assign _T_11096 = 5'he == _T_10211_20; // @[Mux.scala 46:19:@9760.4]
  assign _T_11097 = _T_11096 ? _T_9260_13 : _T_11095; // @[Mux.scala 46:16:@9761.4]
  assign _T_11098 = 5'hd == _T_10211_20; // @[Mux.scala 46:19:@9762.4]
  assign _T_11099 = _T_11098 ? _T_9260_12 : _T_11097; // @[Mux.scala 46:16:@9763.4]
  assign _T_11100 = 5'hc == _T_10211_20; // @[Mux.scala 46:19:@9764.4]
  assign _T_11101 = _T_11100 ? _T_9260_11 : _T_11099; // @[Mux.scala 46:16:@9765.4]
  assign _T_11102 = 5'hb == _T_10211_20; // @[Mux.scala 46:19:@9766.4]
  assign _T_11103 = _T_11102 ? _T_9260_10 : _T_11101; // @[Mux.scala 46:16:@9767.4]
  assign _T_11104 = 5'ha == _T_10211_20; // @[Mux.scala 46:19:@9768.4]
  assign _T_11105 = _T_11104 ? _T_9260_9 : _T_11103; // @[Mux.scala 46:16:@9769.4]
  assign _T_11106 = 5'h9 == _T_10211_20; // @[Mux.scala 46:19:@9770.4]
  assign _T_11107 = _T_11106 ? _T_9260_8 : _T_11105; // @[Mux.scala 46:16:@9771.4]
  assign _T_11108 = 5'h8 == _T_10211_20; // @[Mux.scala 46:19:@9772.4]
  assign _T_11109 = _T_11108 ? _T_9260_7 : _T_11107; // @[Mux.scala 46:16:@9773.4]
  assign _T_11110 = 5'h7 == _T_10211_20; // @[Mux.scala 46:19:@9774.4]
  assign _T_11111 = _T_11110 ? _T_9260_6 : _T_11109; // @[Mux.scala 46:16:@9775.4]
  assign _T_11112 = 5'h6 == _T_10211_20; // @[Mux.scala 46:19:@9776.4]
  assign _T_11113 = _T_11112 ? _T_9260_5 : _T_11111; // @[Mux.scala 46:16:@9777.4]
  assign _T_11114 = 5'h5 == _T_10211_20; // @[Mux.scala 46:19:@9778.4]
  assign _T_11115 = _T_11114 ? _T_9260_4 : _T_11113; // @[Mux.scala 46:16:@9779.4]
  assign _T_11116 = 5'h4 == _T_10211_20; // @[Mux.scala 46:19:@9780.4]
  assign _T_11117 = _T_11116 ? _T_9260_3 : _T_11115; // @[Mux.scala 46:16:@9781.4]
  assign _T_11118 = 5'h3 == _T_10211_20; // @[Mux.scala 46:19:@9782.4]
  assign _T_11119 = _T_11118 ? _T_9260_2 : _T_11117; // @[Mux.scala 46:16:@9783.4]
  assign _T_11120 = 5'h2 == _T_10211_20; // @[Mux.scala 46:19:@9784.4]
  assign _T_11121 = _T_11120 ? _T_9260_1 : _T_11119; // @[Mux.scala 46:16:@9785.4]
  assign _T_11122 = 5'h1 == _T_10211_20; // @[Mux.scala 46:19:@9786.4]
  assign _T_11123 = _T_11122 ? _T_9260_0 : _T_11121; // @[Mux.scala 46:16:@9787.4]
  assign _T_11147 = 5'h16 == _T_10211_21; // @[Mux.scala 46:19:@9789.4]
  assign _T_11148 = _T_11147 ? _T_9260_21 : 8'h0; // @[Mux.scala 46:16:@9790.4]
  assign _T_11149 = 5'h15 == _T_10211_21; // @[Mux.scala 46:19:@9791.4]
  assign _T_11150 = _T_11149 ? _T_9260_20 : _T_11148; // @[Mux.scala 46:16:@9792.4]
  assign _T_11151 = 5'h14 == _T_10211_21; // @[Mux.scala 46:19:@9793.4]
  assign _T_11152 = _T_11151 ? _T_9260_19 : _T_11150; // @[Mux.scala 46:16:@9794.4]
  assign _T_11153 = 5'h13 == _T_10211_21; // @[Mux.scala 46:19:@9795.4]
  assign _T_11154 = _T_11153 ? _T_9260_18 : _T_11152; // @[Mux.scala 46:16:@9796.4]
  assign _T_11155 = 5'h12 == _T_10211_21; // @[Mux.scala 46:19:@9797.4]
  assign _T_11156 = _T_11155 ? _T_9260_17 : _T_11154; // @[Mux.scala 46:16:@9798.4]
  assign _T_11157 = 5'h11 == _T_10211_21; // @[Mux.scala 46:19:@9799.4]
  assign _T_11158 = _T_11157 ? _T_9260_16 : _T_11156; // @[Mux.scala 46:16:@9800.4]
  assign _T_11159 = 5'h10 == _T_10211_21; // @[Mux.scala 46:19:@9801.4]
  assign _T_11160 = _T_11159 ? _T_9260_15 : _T_11158; // @[Mux.scala 46:16:@9802.4]
  assign _T_11161 = 5'hf == _T_10211_21; // @[Mux.scala 46:19:@9803.4]
  assign _T_11162 = _T_11161 ? _T_9260_14 : _T_11160; // @[Mux.scala 46:16:@9804.4]
  assign _T_11163 = 5'he == _T_10211_21; // @[Mux.scala 46:19:@9805.4]
  assign _T_11164 = _T_11163 ? _T_9260_13 : _T_11162; // @[Mux.scala 46:16:@9806.4]
  assign _T_11165 = 5'hd == _T_10211_21; // @[Mux.scala 46:19:@9807.4]
  assign _T_11166 = _T_11165 ? _T_9260_12 : _T_11164; // @[Mux.scala 46:16:@9808.4]
  assign _T_11167 = 5'hc == _T_10211_21; // @[Mux.scala 46:19:@9809.4]
  assign _T_11168 = _T_11167 ? _T_9260_11 : _T_11166; // @[Mux.scala 46:16:@9810.4]
  assign _T_11169 = 5'hb == _T_10211_21; // @[Mux.scala 46:19:@9811.4]
  assign _T_11170 = _T_11169 ? _T_9260_10 : _T_11168; // @[Mux.scala 46:16:@9812.4]
  assign _T_11171 = 5'ha == _T_10211_21; // @[Mux.scala 46:19:@9813.4]
  assign _T_11172 = _T_11171 ? _T_9260_9 : _T_11170; // @[Mux.scala 46:16:@9814.4]
  assign _T_11173 = 5'h9 == _T_10211_21; // @[Mux.scala 46:19:@9815.4]
  assign _T_11174 = _T_11173 ? _T_9260_8 : _T_11172; // @[Mux.scala 46:16:@9816.4]
  assign _T_11175 = 5'h8 == _T_10211_21; // @[Mux.scala 46:19:@9817.4]
  assign _T_11176 = _T_11175 ? _T_9260_7 : _T_11174; // @[Mux.scala 46:16:@9818.4]
  assign _T_11177 = 5'h7 == _T_10211_21; // @[Mux.scala 46:19:@9819.4]
  assign _T_11178 = _T_11177 ? _T_9260_6 : _T_11176; // @[Mux.scala 46:16:@9820.4]
  assign _T_11179 = 5'h6 == _T_10211_21; // @[Mux.scala 46:19:@9821.4]
  assign _T_11180 = _T_11179 ? _T_9260_5 : _T_11178; // @[Mux.scala 46:16:@9822.4]
  assign _T_11181 = 5'h5 == _T_10211_21; // @[Mux.scala 46:19:@9823.4]
  assign _T_11182 = _T_11181 ? _T_9260_4 : _T_11180; // @[Mux.scala 46:16:@9824.4]
  assign _T_11183 = 5'h4 == _T_10211_21; // @[Mux.scala 46:19:@9825.4]
  assign _T_11184 = _T_11183 ? _T_9260_3 : _T_11182; // @[Mux.scala 46:16:@9826.4]
  assign _T_11185 = 5'h3 == _T_10211_21; // @[Mux.scala 46:19:@9827.4]
  assign _T_11186 = _T_11185 ? _T_9260_2 : _T_11184; // @[Mux.scala 46:16:@9828.4]
  assign _T_11187 = 5'h2 == _T_10211_21; // @[Mux.scala 46:19:@9829.4]
  assign _T_11188 = _T_11187 ? _T_9260_1 : _T_11186; // @[Mux.scala 46:16:@9830.4]
  assign _T_11189 = 5'h1 == _T_10211_21; // @[Mux.scala 46:19:@9831.4]
  assign _T_11190 = _T_11189 ? _T_9260_0 : _T_11188; // @[Mux.scala 46:16:@9832.4]
  assign _T_11215 = 5'h17 == _T_10211_22; // @[Mux.scala 46:19:@9834.4]
  assign _T_11216 = _T_11215 ? _T_9260_22 : 8'h0; // @[Mux.scala 46:16:@9835.4]
  assign _T_11217 = 5'h16 == _T_10211_22; // @[Mux.scala 46:19:@9836.4]
  assign _T_11218 = _T_11217 ? _T_9260_21 : _T_11216; // @[Mux.scala 46:16:@9837.4]
  assign _T_11219 = 5'h15 == _T_10211_22; // @[Mux.scala 46:19:@9838.4]
  assign _T_11220 = _T_11219 ? _T_9260_20 : _T_11218; // @[Mux.scala 46:16:@9839.4]
  assign _T_11221 = 5'h14 == _T_10211_22; // @[Mux.scala 46:19:@9840.4]
  assign _T_11222 = _T_11221 ? _T_9260_19 : _T_11220; // @[Mux.scala 46:16:@9841.4]
  assign _T_11223 = 5'h13 == _T_10211_22; // @[Mux.scala 46:19:@9842.4]
  assign _T_11224 = _T_11223 ? _T_9260_18 : _T_11222; // @[Mux.scala 46:16:@9843.4]
  assign _T_11225 = 5'h12 == _T_10211_22; // @[Mux.scala 46:19:@9844.4]
  assign _T_11226 = _T_11225 ? _T_9260_17 : _T_11224; // @[Mux.scala 46:16:@9845.4]
  assign _T_11227 = 5'h11 == _T_10211_22; // @[Mux.scala 46:19:@9846.4]
  assign _T_11228 = _T_11227 ? _T_9260_16 : _T_11226; // @[Mux.scala 46:16:@9847.4]
  assign _T_11229 = 5'h10 == _T_10211_22; // @[Mux.scala 46:19:@9848.4]
  assign _T_11230 = _T_11229 ? _T_9260_15 : _T_11228; // @[Mux.scala 46:16:@9849.4]
  assign _T_11231 = 5'hf == _T_10211_22; // @[Mux.scala 46:19:@9850.4]
  assign _T_11232 = _T_11231 ? _T_9260_14 : _T_11230; // @[Mux.scala 46:16:@9851.4]
  assign _T_11233 = 5'he == _T_10211_22; // @[Mux.scala 46:19:@9852.4]
  assign _T_11234 = _T_11233 ? _T_9260_13 : _T_11232; // @[Mux.scala 46:16:@9853.4]
  assign _T_11235 = 5'hd == _T_10211_22; // @[Mux.scala 46:19:@9854.4]
  assign _T_11236 = _T_11235 ? _T_9260_12 : _T_11234; // @[Mux.scala 46:16:@9855.4]
  assign _T_11237 = 5'hc == _T_10211_22; // @[Mux.scala 46:19:@9856.4]
  assign _T_11238 = _T_11237 ? _T_9260_11 : _T_11236; // @[Mux.scala 46:16:@9857.4]
  assign _T_11239 = 5'hb == _T_10211_22; // @[Mux.scala 46:19:@9858.4]
  assign _T_11240 = _T_11239 ? _T_9260_10 : _T_11238; // @[Mux.scala 46:16:@9859.4]
  assign _T_11241 = 5'ha == _T_10211_22; // @[Mux.scala 46:19:@9860.4]
  assign _T_11242 = _T_11241 ? _T_9260_9 : _T_11240; // @[Mux.scala 46:16:@9861.4]
  assign _T_11243 = 5'h9 == _T_10211_22; // @[Mux.scala 46:19:@9862.4]
  assign _T_11244 = _T_11243 ? _T_9260_8 : _T_11242; // @[Mux.scala 46:16:@9863.4]
  assign _T_11245 = 5'h8 == _T_10211_22; // @[Mux.scala 46:19:@9864.4]
  assign _T_11246 = _T_11245 ? _T_9260_7 : _T_11244; // @[Mux.scala 46:16:@9865.4]
  assign _T_11247 = 5'h7 == _T_10211_22; // @[Mux.scala 46:19:@9866.4]
  assign _T_11248 = _T_11247 ? _T_9260_6 : _T_11246; // @[Mux.scala 46:16:@9867.4]
  assign _T_11249 = 5'h6 == _T_10211_22; // @[Mux.scala 46:19:@9868.4]
  assign _T_11250 = _T_11249 ? _T_9260_5 : _T_11248; // @[Mux.scala 46:16:@9869.4]
  assign _T_11251 = 5'h5 == _T_10211_22; // @[Mux.scala 46:19:@9870.4]
  assign _T_11252 = _T_11251 ? _T_9260_4 : _T_11250; // @[Mux.scala 46:16:@9871.4]
  assign _T_11253 = 5'h4 == _T_10211_22; // @[Mux.scala 46:19:@9872.4]
  assign _T_11254 = _T_11253 ? _T_9260_3 : _T_11252; // @[Mux.scala 46:16:@9873.4]
  assign _T_11255 = 5'h3 == _T_10211_22; // @[Mux.scala 46:19:@9874.4]
  assign _T_11256 = _T_11255 ? _T_9260_2 : _T_11254; // @[Mux.scala 46:16:@9875.4]
  assign _T_11257 = 5'h2 == _T_10211_22; // @[Mux.scala 46:19:@9876.4]
  assign _T_11258 = _T_11257 ? _T_9260_1 : _T_11256; // @[Mux.scala 46:16:@9877.4]
  assign _T_11259 = 5'h1 == _T_10211_22; // @[Mux.scala 46:19:@9878.4]
  assign _T_11260 = _T_11259 ? _T_9260_0 : _T_11258; // @[Mux.scala 46:16:@9879.4]
  assign _T_11286 = 5'h18 == _T_10211_23; // @[Mux.scala 46:19:@9881.4]
  assign _T_11287 = _T_11286 ? _T_9260_23 : 8'h0; // @[Mux.scala 46:16:@9882.4]
  assign _T_11288 = 5'h17 == _T_10211_23; // @[Mux.scala 46:19:@9883.4]
  assign _T_11289 = _T_11288 ? _T_9260_22 : _T_11287; // @[Mux.scala 46:16:@9884.4]
  assign _T_11290 = 5'h16 == _T_10211_23; // @[Mux.scala 46:19:@9885.4]
  assign _T_11291 = _T_11290 ? _T_9260_21 : _T_11289; // @[Mux.scala 46:16:@9886.4]
  assign _T_11292 = 5'h15 == _T_10211_23; // @[Mux.scala 46:19:@9887.4]
  assign _T_11293 = _T_11292 ? _T_9260_20 : _T_11291; // @[Mux.scala 46:16:@9888.4]
  assign _T_11294 = 5'h14 == _T_10211_23; // @[Mux.scala 46:19:@9889.4]
  assign _T_11295 = _T_11294 ? _T_9260_19 : _T_11293; // @[Mux.scala 46:16:@9890.4]
  assign _T_11296 = 5'h13 == _T_10211_23; // @[Mux.scala 46:19:@9891.4]
  assign _T_11297 = _T_11296 ? _T_9260_18 : _T_11295; // @[Mux.scala 46:16:@9892.4]
  assign _T_11298 = 5'h12 == _T_10211_23; // @[Mux.scala 46:19:@9893.4]
  assign _T_11299 = _T_11298 ? _T_9260_17 : _T_11297; // @[Mux.scala 46:16:@9894.4]
  assign _T_11300 = 5'h11 == _T_10211_23; // @[Mux.scala 46:19:@9895.4]
  assign _T_11301 = _T_11300 ? _T_9260_16 : _T_11299; // @[Mux.scala 46:16:@9896.4]
  assign _T_11302 = 5'h10 == _T_10211_23; // @[Mux.scala 46:19:@9897.4]
  assign _T_11303 = _T_11302 ? _T_9260_15 : _T_11301; // @[Mux.scala 46:16:@9898.4]
  assign _T_11304 = 5'hf == _T_10211_23; // @[Mux.scala 46:19:@9899.4]
  assign _T_11305 = _T_11304 ? _T_9260_14 : _T_11303; // @[Mux.scala 46:16:@9900.4]
  assign _T_11306 = 5'he == _T_10211_23; // @[Mux.scala 46:19:@9901.4]
  assign _T_11307 = _T_11306 ? _T_9260_13 : _T_11305; // @[Mux.scala 46:16:@9902.4]
  assign _T_11308 = 5'hd == _T_10211_23; // @[Mux.scala 46:19:@9903.4]
  assign _T_11309 = _T_11308 ? _T_9260_12 : _T_11307; // @[Mux.scala 46:16:@9904.4]
  assign _T_11310 = 5'hc == _T_10211_23; // @[Mux.scala 46:19:@9905.4]
  assign _T_11311 = _T_11310 ? _T_9260_11 : _T_11309; // @[Mux.scala 46:16:@9906.4]
  assign _T_11312 = 5'hb == _T_10211_23; // @[Mux.scala 46:19:@9907.4]
  assign _T_11313 = _T_11312 ? _T_9260_10 : _T_11311; // @[Mux.scala 46:16:@9908.4]
  assign _T_11314 = 5'ha == _T_10211_23; // @[Mux.scala 46:19:@9909.4]
  assign _T_11315 = _T_11314 ? _T_9260_9 : _T_11313; // @[Mux.scala 46:16:@9910.4]
  assign _T_11316 = 5'h9 == _T_10211_23; // @[Mux.scala 46:19:@9911.4]
  assign _T_11317 = _T_11316 ? _T_9260_8 : _T_11315; // @[Mux.scala 46:16:@9912.4]
  assign _T_11318 = 5'h8 == _T_10211_23; // @[Mux.scala 46:19:@9913.4]
  assign _T_11319 = _T_11318 ? _T_9260_7 : _T_11317; // @[Mux.scala 46:16:@9914.4]
  assign _T_11320 = 5'h7 == _T_10211_23; // @[Mux.scala 46:19:@9915.4]
  assign _T_11321 = _T_11320 ? _T_9260_6 : _T_11319; // @[Mux.scala 46:16:@9916.4]
  assign _T_11322 = 5'h6 == _T_10211_23; // @[Mux.scala 46:19:@9917.4]
  assign _T_11323 = _T_11322 ? _T_9260_5 : _T_11321; // @[Mux.scala 46:16:@9918.4]
  assign _T_11324 = 5'h5 == _T_10211_23; // @[Mux.scala 46:19:@9919.4]
  assign _T_11325 = _T_11324 ? _T_9260_4 : _T_11323; // @[Mux.scala 46:16:@9920.4]
  assign _T_11326 = 5'h4 == _T_10211_23; // @[Mux.scala 46:19:@9921.4]
  assign _T_11327 = _T_11326 ? _T_9260_3 : _T_11325; // @[Mux.scala 46:16:@9922.4]
  assign _T_11328 = 5'h3 == _T_10211_23; // @[Mux.scala 46:19:@9923.4]
  assign _T_11329 = _T_11328 ? _T_9260_2 : _T_11327; // @[Mux.scala 46:16:@9924.4]
  assign _T_11330 = 5'h2 == _T_10211_23; // @[Mux.scala 46:19:@9925.4]
  assign _T_11331 = _T_11330 ? _T_9260_1 : _T_11329; // @[Mux.scala 46:16:@9926.4]
  assign _T_11332 = 5'h1 == _T_10211_23; // @[Mux.scala 46:19:@9927.4]
  assign _T_11333 = _T_11332 ? _T_9260_0 : _T_11331; // @[Mux.scala 46:16:@9928.4]
  assign _T_11360 = 5'h19 == _T_10211_24; // @[Mux.scala 46:19:@9930.4]
  assign _T_11361 = _T_11360 ? _T_9260_24 : 8'h0; // @[Mux.scala 46:16:@9931.4]
  assign _T_11362 = 5'h18 == _T_10211_24; // @[Mux.scala 46:19:@9932.4]
  assign _T_11363 = _T_11362 ? _T_9260_23 : _T_11361; // @[Mux.scala 46:16:@9933.4]
  assign _T_11364 = 5'h17 == _T_10211_24; // @[Mux.scala 46:19:@9934.4]
  assign _T_11365 = _T_11364 ? _T_9260_22 : _T_11363; // @[Mux.scala 46:16:@9935.4]
  assign _T_11366 = 5'h16 == _T_10211_24; // @[Mux.scala 46:19:@9936.4]
  assign _T_11367 = _T_11366 ? _T_9260_21 : _T_11365; // @[Mux.scala 46:16:@9937.4]
  assign _T_11368 = 5'h15 == _T_10211_24; // @[Mux.scala 46:19:@9938.4]
  assign _T_11369 = _T_11368 ? _T_9260_20 : _T_11367; // @[Mux.scala 46:16:@9939.4]
  assign _T_11370 = 5'h14 == _T_10211_24; // @[Mux.scala 46:19:@9940.4]
  assign _T_11371 = _T_11370 ? _T_9260_19 : _T_11369; // @[Mux.scala 46:16:@9941.4]
  assign _T_11372 = 5'h13 == _T_10211_24; // @[Mux.scala 46:19:@9942.4]
  assign _T_11373 = _T_11372 ? _T_9260_18 : _T_11371; // @[Mux.scala 46:16:@9943.4]
  assign _T_11374 = 5'h12 == _T_10211_24; // @[Mux.scala 46:19:@9944.4]
  assign _T_11375 = _T_11374 ? _T_9260_17 : _T_11373; // @[Mux.scala 46:16:@9945.4]
  assign _T_11376 = 5'h11 == _T_10211_24; // @[Mux.scala 46:19:@9946.4]
  assign _T_11377 = _T_11376 ? _T_9260_16 : _T_11375; // @[Mux.scala 46:16:@9947.4]
  assign _T_11378 = 5'h10 == _T_10211_24; // @[Mux.scala 46:19:@9948.4]
  assign _T_11379 = _T_11378 ? _T_9260_15 : _T_11377; // @[Mux.scala 46:16:@9949.4]
  assign _T_11380 = 5'hf == _T_10211_24; // @[Mux.scala 46:19:@9950.4]
  assign _T_11381 = _T_11380 ? _T_9260_14 : _T_11379; // @[Mux.scala 46:16:@9951.4]
  assign _T_11382 = 5'he == _T_10211_24; // @[Mux.scala 46:19:@9952.4]
  assign _T_11383 = _T_11382 ? _T_9260_13 : _T_11381; // @[Mux.scala 46:16:@9953.4]
  assign _T_11384 = 5'hd == _T_10211_24; // @[Mux.scala 46:19:@9954.4]
  assign _T_11385 = _T_11384 ? _T_9260_12 : _T_11383; // @[Mux.scala 46:16:@9955.4]
  assign _T_11386 = 5'hc == _T_10211_24; // @[Mux.scala 46:19:@9956.4]
  assign _T_11387 = _T_11386 ? _T_9260_11 : _T_11385; // @[Mux.scala 46:16:@9957.4]
  assign _T_11388 = 5'hb == _T_10211_24; // @[Mux.scala 46:19:@9958.4]
  assign _T_11389 = _T_11388 ? _T_9260_10 : _T_11387; // @[Mux.scala 46:16:@9959.4]
  assign _T_11390 = 5'ha == _T_10211_24; // @[Mux.scala 46:19:@9960.4]
  assign _T_11391 = _T_11390 ? _T_9260_9 : _T_11389; // @[Mux.scala 46:16:@9961.4]
  assign _T_11392 = 5'h9 == _T_10211_24; // @[Mux.scala 46:19:@9962.4]
  assign _T_11393 = _T_11392 ? _T_9260_8 : _T_11391; // @[Mux.scala 46:16:@9963.4]
  assign _T_11394 = 5'h8 == _T_10211_24; // @[Mux.scala 46:19:@9964.4]
  assign _T_11395 = _T_11394 ? _T_9260_7 : _T_11393; // @[Mux.scala 46:16:@9965.4]
  assign _T_11396 = 5'h7 == _T_10211_24; // @[Mux.scala 46:19:@9966.4]
  assign _T_11397 = _T_11396 ? _T_9260_6 : _T_11395; // @[Mux.scala 46:16:@9967.4]
  assign _T_11398 = 5'h6 == _T_10211_24; // @[Mux.scala 46:19:@9968.4]
  assign _T_11399 = _T_11398 ? _T_9260_5 : _T_11397; // @[Mux.scala 46:16:@9969.4]
  assign _T_11400 = 5'h5 == _T_10211_24; // @[Mux.scala 46:19:@9970.4]
  assign _T_11401 = _T_11400 ? _T_9260_4 : _T_11399; // @[Mux.scala 46:16:@9971.4]
  assign _T_11402 = 5'h4 == _T_10211_24; // @[Mux.scala 46:19:@9972.4]
  assign _T_11403 = _T_11402 ? _T_9260_3 : _T_11401; // @[Mux.scala 46:16:@9973.4]
  assign _T_11404 = 5'h3 == _T_10211_24; // @[Mux.scala 46:19:@9974.4]
  assign _T_11405 = _T_11404 ? _T_9260_2 : _T_11403; // @[Mux.scala 46:16:@9975.4]
  assign _T_11406 = 5'h2 == _T_10211_24; // @[Mux.scala 46:19:@9976.4]
  assign _T_11407 = _T_11406 ? _T_9260_1 : _T_11405; // @[Mux.scala 46:16:@9977.4]
  assign _T_11408 = 5'h1 == _T_10211_24; // @[Mux.scala 46:19:@9978.4]
  assign _T_11409 = _T_11408 ? _T_9260_0 : _T_11407; // @[Mux.scala 46:16:@9979.4]
  assign _T_11437 = 5'h1a == _T_10211_25; // @[Mux.scala 46:19:@9981.4]
  assign _T_11438 = _T_11437 ? _T_9260_25 : 8'h0; // @[Mux.scala 46:16:@9982.4]
  assign _T_11439 = 5'h19 == _T_10211_25; // @[Mux.scala 46:19:@9983.4]
  assign _T_11440 = _T_11439 ? _T_9260_24 : _T_11438; // @[Mux.scala 46:16:@9984.4]
  assign _T_11441 = 5'h18 == _T_10211_25; // @[Mux.scala 46:19:@9985.4]
  assign _T_11442 = _T_11441 ? _T_9260_23 : _T_11440; // @[Mux.scala 46:16:@9986.4]
  assign _T_11443 = 5'h17 == _T_10211_25; // @[Mux.scala 46:19:@9987.4]
  assign _T_11444 = _T_11443 ? _T_9260_22 : _T_11442; // @[Mux.scala 46:16:@9988.4]
  assign _T_11445 = 5'h16 == _T_10211_25; // @[Mux.scala 46:19:@9989.4]
  assign _T_11446 = _T_11445 ? _T_9260_21 : _T_11444; // @[Mux.scala 46:16:@9990.4]
  assign _T_11447 = 5'h15 == _T_10211_25; // @[Mux.scala 46:19:@9991.4]
  assign _T_11448 = _T_11447 ? _T_9260_20 : _T_11446; // @[Mux.scala 46:16:@9992.4]
  assign _T_11449 = 5'h14 == _T_10211_25; // @[Mux.scala 46:19:@9993.4]
  assign _T_11450 = _T_11449 ? _T_9260_19 : _T_11448; // @[Mux.scala 46:16:@9994.4]
  assign _T_11451 = 5'h13 == _T_10211_25; // @[Mux.scala 46:19:@9995.4]
  assign _T_11452 = _T_11451 ? _T_9260_18 : _T_11450; // @[Mux.scala 46:16:@9996.4]
  assign _T_11453 = 5'h12 == _T_10211_25; // @[Mux.scala 46:19:@9997.4]
  assign _T_11454 = _T_11453 ? _T_9260_17 : _T_11452; // @[Mux.scala 46:16:@9998.4]
  assign _T_11455 = 5'h11 == _T_10211_25; // @[Mux.scala 46:19:@9999.4]
  assign _T_11456 = _T_11455 ? _T_9260_16 : _T_11454; // @[Mux.scala 46:16:@10000.4]
  assign _T_11457 = 5'h10 == _T_10211_25; // @[Mux.scala 46:19:@10001.4]
  assign _T_11458 = _T_11457 ? _T_9260_15 : _T_11456; // @[Mux.scala 46:16:@10002.4]
  assign _T_11459 = 5'hf == _T_10211_25; // @[Mux.scala 46:19:@10003.4]
  assign _T_11460 = _T_11459 ? _T_9260_14 : _T_11458; // @[Mux.scala 46:16:@10004.4]
  assign _T_11461 = 5'he == _T_10211_25; // @[Mux.scala 46:19:@10005.4]
  assign _T_11462 = _T_11461 ? _T_9260_13 : _T_11460; // @[Mux.scala 46:16:@10006.4]
  assign _T_11463 = 5'hd == _T_10211_25; // @[Mux.scala 46:19:@10007.4]
  assign _T_11464 = _T_11463 ? _T_9260_12 : _T_11462; // @[Mux.scala 46:16:@10008.4]
  assign _T_11465 = 5'hc == _T_10211_25; // @[Mux.scala 46:19:@10009.4]
  assign _T_11466 = _T_11465 ? _T_9260_11 : _T_11464; // @[Mux.scala 46:16:@10010.4]
  assign _T_11467 = 5'hb == _T_10211_25; // @[Mux.scala 46:19:@10011.4]
  assign _T_11468 = _T_11467 ? _T_9260_10 : _T_11466; // @[Mux.scala 46:16:@10012.4]
  assign _T_11469 = 5'ha == _T_10211_25; // @[Mux.scala 46:19:@10013.4]
  assign _T_11470 = _T_11469 ? _T_9260_9 : _T_11468; // @[Mux.scala 46:16:@10014.4]
  assign _T_11471 = 5'h9 == _T_10211_25; // @[Mux.scala 46:19:@10015.4]
  assign _T_11472 = _T_11471 ? _T_9260_8 : _T_11470; // @[Mux.scala 46:16:@10016.4]
  assign _T_11473 = 5'h8 == _T_10211_25; // @[Mux.scala 46:19:@10017.4]
  assign _T_11474 = _T_11473 ? _T_9260_7 : _T_11472; // @[Mux.scala 46:16:@10018.4]
  assign _T_11475 = 5'h7 == _T_10211_25; // @[Mux.scala 46:19:@10019.4]
  assign _T_11476 = _T_11475 ? _T_9260_6 : _T_11474; // @[Mux.scala 46:16:@10020.4]
  assign _T_11477 = 5'h6 == _T_10211_25; // @[Mux.scala 46:19:@10021.4]
  assign _T_11478 = _T_11477 ? _T_9260_5 : _T_11476; // @[Mux.scala 46:16:@10022.4]
  assign _T_11479 = 5'h5 == _T_10211_25; // @[Mux.scala 46:19:@10023.4]
  assign _T_11480 = _T_11479 ? _T_9260_4 : _T_11478; // @[Mux.scala 46:16:@10024.4]
  assign _T_11481 = 5'h4 == _T_10211_25; // @[Mux.scala 46:19:@10025.4]
  assign _T_11482 = _T_11481 ? _T_9260_3 : _T_11480; // @[Mux.scala 46:16:@10026.4]
  assign _T_11483 = 5'h3 == _T_10211_25; // @[Mux.scala 46:19:@10027.4]
  assign _T_11484 = _T_11483 ? _T_9260_2 : _T_11482; // @[Mux.scala 46:16:@10028.4]
  assign _T_11485 = 5'h2 == _T_10211_25; // @[Mux.scala 46:19:@10029.4]
  assign _T_11486 = _T_11485 ? _T_9260_1 : _T_11484; // @[Mux.scala 46:16:@10030.4]
  assign _T_11487 = 5'h1 == _T_10211_25; // @[Mux.scala 46:19:@10031.4]
  assign _T_11488 = _T_11487 ? _T_9260_0 : _T_11486; // @[Mux.scala 46:16:@10032.4]
  assign _T_11517 = 5'h1b == _T_10211_26; // @[Mux.scala 46:19:@10034.4]
  assign _T_11518 = _T_11517 ? _T_9260_26 : 8'h0; // @[Mux.scala 46:16:@10035.4]
  assign _T_11519 = 5'h1a == _T_10211_26; // @[Mux.scala 46:19:@10036.4]
  assign _T_11520 = _T_11519 ? _T_9260_25 : _T_11518; // @[Mux.scala 46:16:@10037.4]
  assign _T_11521 = 5'h19 == _T_10211_26; // @[Mux.scala 46:19:@10038.4]
  assign _T_11522 = _T_11521 ? _T_9260_24 : _T_11520; // @[Mux.scala 46:16:@10039.4]
  assign _T_11523 = 5'h18 == _T_10211_26; // @[Mux.scala 46:19:@10040.4]
  assign _T_11524 = _T_11523 ? _T_9260_23 : _T_11522; // @[Mux.scala 46:16:@10041.4]
  assign _T_11525 = 5'h17 == _T_10211_26; // @[Mux.scala 46:19:@10042.4]
  assign _T_11526 = _T_11525 ? _T_9260_22 : _T_11524; // @[Mux.scala 46:16:@10043.4]
  assign _T_11527 = 5'h16 == _T_10211_26; // @[Mux.scala 46:19:@10044.4]
  assign _T_11528 = _T_11527 ? _T_9260_21 : _T_11526; // @[Mux.scala 46:16:@10045.4]
  assign _T_11529 = 5'h15 == _T_10211_26; // @[Mux.scala 46:19:@10046.4]
  assign _T_11530 = _T_11529 ? _T_9260_20 : _T_11528; // @[Mux.scala 46:16:@10047.4]
  assign _T_11531 = 5'h14 == _T_10211_26; // @[Mux.scala 46:19:@10048.4]
  assign _T_11532 = _T_11531 ? _T_9260_19 : _T_11530; // @[Mux.scala 46:16:@10049.4]
  assign _T_11533 = 5'h13 == _T_10211_26; // @[Mux.scala 46:19:@10050.4]
  assign _T_11534 = _T_11533 ? _T_9260_18 : _T_11532; // @[Mux.scala 46:16:@10051.4]
  assign _T_11535 = 5'h12 == _T_10211_26; // @[Mux.scala 46:19:@10052.4]
  assign _T_11536 = _T_11535 ? _T_9260_17 : _T_11534; // @[Mux.scala 46:16:@10053.4]
  assign _T_11537 = 5'h11 == _T_10211_26; // @[Mux.scala 46:19:@10054.4]
  assign _T_11538 = _T_11537 ? _T_9260_16 : _T_11536; // @[Mux.scala 46:16:@10055.4]
  assign _T_11539 = 5'h10 == _T_10211_26; // @[Mux.scala 46:19:@10056.4]
  assign _T_11540 = _T_11539 ? _T_9260_15 : _T_11538; // @[Mux.scala 46:16:@10057.4]
  assign _T_11541 = 5'hf == _T_10211_26; // @[Mux.scala 46:19:@10058.4]
  assign _T_11542 = _T_11541 ? _T_9260_14 : _T_11540; // @[Mux.scala 46:16:@10059.4]
  assign _T_11543 = 5'he == _T_10211_26; // @[Mux.scala 46:19:@10060.4]
  assign _T_11544 = _T_11543 ? _T_9260_13 : _T_11542; // @[Mux.scala 46:16:@10061.4]
  assign _T_11545 = 5'hd == _T_10211_26; // @[Mux.scala 46:19:@10062.4]
  assign _T_11546 = _T_11545 ? _T_9260_12 : _T_11544; // @[Mux.scala 46:16:@10063.4]
  assign _T_11547 = 5'hc == _T_10211_26; // @[Mux.scala 46:19:@10064.4]
  assign _T_11548 = _T_11547 ? _T_9260_11 : _T_11546; // @[Mux.scala 46:16:@10065.4]
  assign _T_11549 = 5'hb == _T_10211_26; // @[Mux.scala 46:19:@10066.4]
  assign _T_11550 = _T_11549 ? _T_9260_10 : _T_11548; // @[Mux.scala 46:16:@10067.4]
  assign _T_11551 = 5'ha == _T_10211_26; // @[Mux.scala 46:19:@10068.4]
  assign _T_11552 = _T_11551 ? _T_9260_9 : _T_11550; // @[Mux.scala 46:16:@10069.4]
  assign _T_11553 = 5'h9 == _T_10211_26; // @[Mux.scala 46:19:@10070.4]
  assign _T_11554 = _T_11553 ? _T_9260_8 : _T_11552; // @[Mux.scala 46:16:@10071.4]
  assign _T_11555 = 5'h8 == _T_10211_26; // @[Mux.scala 46:19:@10072.4]
  assign _T_11556 = _T_11555 ? _T_9260_7 : _T_11554; // @[Mux.scala 46:16:@10073.4]
  assign _T_11557 = 5'h7 == _T_10211_26; // @[Mux.scala 46:19:@10074.4]
  assign _T_11558 = _T_11557 ? _T_9260_6 : _T_11556; // @[Mux.scala 46:16:@10075.4]
  assign _T_11559 = 5'h6 == _T_10211_26; // @[Mux.scala 46:19:@10076.4]
  assign _T_11560 = _T_11559 ? _T_9260_5 : _T_11558; // @[Mux.scala 46:16:@10077.4]
  assign _T_11561 = 5'h5 == _T_10211_26; // @[Mux.scala 46:19:@10078.4]
  assign _T_11562 = _T_11561 ? _T_9260_4 : _T_11560; // @[Mux.scala 46:16:@10079.4]
  assign _T_11563 = 5'h4 == _T_10211_26; // @[Mux.scala 46:19:@10080.4]
  assign _T_11564 = _T_11563 ? _T_9260_3 : _T_11562; // @[Mux.scala 46:16:@10081.4]
  assign _T_11565 = 5'h3 == _T_10211_26; // @[Mux.scala 46:19:@10082.4]
  assign _T_11566 = _T_11565 ? _T_9260_2 : _T_11564; // @[Mux.scala 46:16:@10083.4]
  assign _T_11567 = 5'h2 == _T_10211_26; // @[Mux.scala 46:19:@10084.4]
  assign _T_11568 = _T_11567 ? _T_9260_1 : _T_11566; // @[Mux.scala 46:16:@10085.4]
  assign _T_11569 = 5'h1 == _T_10211_26; // @[Mux.scala 46:19:@10086.4]
  assign _T_11570 = _T_11569 ? _T_9260_0 : _T_11568; // @[Mux.scala 46:16:@10087.4]
  assign _T_11600 = 5'h1c == _T_10211_27; // @[Mux.scala 46:19:@10089.4]
  assign _T_11601 = _T_11600 ? _T_9260_27 : 8'h0; // @[Mux.scala 46:16:@10090.4]
  assign _T_11602 = 5'h1b == _T_10211_27; // @[Mux.scala 46:19:@10091.4]
  assign _T_11603 = _T_11602 ? _T_9260_26 : _T_11601; // @[Mux.scala 46:16:@10092.4]
  assign _T_11604 = 5'h1a == _T_10211_27; // @[Mux.scala 46:19:@10093.4]
  assign _T_11605 = _T_11604 ? _T_9260_25 : _T_11603; // @[Mux.scala 46:16:@10094.4]
  assign _T_11606 = 5'h19 == _T_10211_27; // @[Mux.scala 46:19:@10095.4]
  assign _T_11607 = _T_11606 ? _T_9260_24 : _T_11605; // @[Mux.scala 46:16:@10096.4]
  assign _T_11608 = 5'h18 == _T_10211_27; // @[Mux.scala 46:19:@10097.4]
  assign _T_11609 = _T_11608 ? _T_9260_23 : _T_11607; // @[Mux.scala 46:16:@10098.4]
  assign _T_11610 = 5'h17 == _T_10211_27; // @[Mux.scala 46:19:@10099.4]
  assign _T_11611 = _T_11610 ? _T_9260_22 : _T_11609; // @[Mux.scala 46:16:@10100.4]
  assign _T_11612 = 5'h16 == _T_10211_27; // @[Mux.scala 46:19:@10101.4]
  assign _T_11613 = _T_11612 ? _T_9260_21 : _T_11611; // @[Mux.scala 46:16:@10102.4]
  assign _T_11614 = 5'h15 == _T_10211_27; // @[Mux.scala 46:19:@10103.4]
  assign _T_11615 = _T_11614 ? _T_9260_20 : _T_11613; // @[Mux.scala 46:16:@10104.4]
  assign _T_11616 = 5'h14 == _T_10211_27; // @[Mux.scala 46:19:@10105.4]
  assign _T_11617 = _T_11616 ? _T_9260_19 : _T_11615; // @[Mux.scala 46:16:@10106.4]
  assign _T_11618 = 5'h13 == _T_10211_27; // @[Mux.scala 46:19:@10107.4]
  assign _T_11619 = _T_11618 ? _T_9260_18 : _T_11617; // @[Mux.scala 46:16:@10108.4]
  assign _T_11620 = 5'h12 == _T_10211_27; // @[Mux.scala 46:19:@10109.4]
  assign _T_11621 = _T_11620 ? _T_9260_17 : _T_11619; // @[Mux.scala 46:16:@10110.4]
  assign _T_11622 = 5'h11 == _T_10211_27; // @[Mux.scala 46:19:@10111.4]
  assign _T_11623 = _T_11622 ? _T_9260_16 : _T_11621; // @[Mux.scala 46:16:@10112.4]
  assign _T_11624 = 5'h10 == _T_10211_27; // @[Mux.scala 46:19:@10113.4]
  assign _T_11625 = _T_11624 ? _T_9260_15 : _T_11623; // @[Mux.scala 46:16:@10114.4]
  assign _T_11626 = 5'hf == _T_10211_27; // @[Mux.scala 46:19:@10115.4]
  assign _T_11627 = _T_11626 ? _T_9260_14 : _T_11625; // @[Mux.scala 46:16:@10116.4]
  assign _T_11628 = 5'he == _T_10211_27; // @[Mux.scala 46:19:@10117.4]
  assign _T_11629 = _T_11628 ? _T_9260_13 : _T_11627; // @[Mux.scala 46:16:@10118.4]
  assign _T_11630 = 5'hd == _T_10211_27; // @[Mux.scala 46:19:@10119.4]
  assign _T_11631 = _T_11630 ? _T_9260_12 : _T_11629; // @[Mux.scala 46:16:@10120.4]
  assign _T_11632 = 5'hc == _T_10211_27; // @[Mux.scala 46:19:@10121.4]
  assign _T_11633 = _T_11632 ? _T_9260_11 : _T_11631; // @[Mux.scala 46:16:@10122.4]
  assign _T_11634 = 5'hb == _T_10211_27; // @[Mux.scala 46:19:@10123.4]
  assign _T_11635 = _T_11634 ? _T_9260_10 : _T_11633; // @[Mux.scala 46:16:@10124.4]
  assign _T_11636 = 5'ha == _T_10211_27; // @[Mux.scala 46:19:@10125.4]
  assign _T_11637 = _T_11636 ? _T_9260_9 : _T_11635; // @[Mux.scala 46:16:@10126.4]
  assign _T_11638 = 5'h9 == _T_10211_27; // @[Mux.scala 46:19:@10127.4]
  assign _T_11639 = _T_11638 ? _T_9260_8 : _T_11637; // @[Mux.scala 46:16:@10128.4]
  assign _T_11640 = 5'h8 == _T_10211_27; // @[Mux.scala 46:19:@10129.4]
  assign _T_11641 = _T_11640 ? _T_9260_7 : _T_11639; // @[Mux.scala 46:16:@10130.4]
  assign _T_11642 = 5'h7 == _T_10211_27; // @[Mux.scala 46:19:@10131.4]
  assign _T_11643 = _T_11642 ? _T_9260_6 : _T_11641; // @[Mux.scala 46:16:@10132.4]
  assign _T_11644 = 5'h6 == _T_10211_27; // @[Mux.scala 46:19:@10133.4]
  assign _T_11645 = _T_11644 ? _T_9260_5 : _T_11643; // @[Mux.scala 46:16:@10134.4]
  assign _T_11646 = 5'h5 == _T_10211_27; // @[Mux.scala 46:19:@10135.4]
  assign _T_11647 = _T_11646 ? _T_9260_4 : _T_11645; // @[Mux.scala 46:16:@10136.4]
  assign _T_11648 = 5'h4 == _T_10211_27; // @[Mux.scala 46:19:@10137.4]
  assign _T_11649 = _T_11648 ? _T_9260_3 : _T_11647; // @[Mux.scala 46:16:@10138.4]
  assign _T_11650 = 5'h3 == _T_10211_27; // @[Mux.scala 46:19:@10139.4]
  assign _T_11651 = _T_11650 ? _T_9260_2 : _T_11649; // @[Mux.scala 46:16:@10140.4]
  assign _T_11652 = 5'h2 == _T_10211_27; // @[Mux.scala 46:19:@10141.4]
  assign _T_11653 = _T_11652 ? _T_9260_1 : _T_11651; // @[Mux.scala 46:16:@10142.4]
  assign _T_11654 = 5'h1 == _T_10211_27; // @[Mux.scala 46:19:@10143.4]
  assign _T_11655 = _T_11654 ? _T_9260_0 : _T_11653; // @[Mux.scala 46:16:@10144.4]
  assign _T_11686 = 5'h1d == _T_10211_28; // @[Mux.scala 46:19:@10146.4]
  assign _T_11687 = _T_11686 ? _T_9260_28 : 8'h0; // @[Mux.scala 46:16:@10147.4]
  assign _T_11688 = 5'h1c == _T_10211_28; // @[Mux.scala 46:19:@10148.4]
  assign _T_11689 = _T_11688 ? _T_9260_27 : _T_11687; // @[Mux.scala 46:16:@10149.4]
  assign _T_11690 = 5'h1b == _T_10211_28; // @[Mux.scala 46:19:@10150.4]
  assign _T_11691 = _T_11690 ? _T_9260_26 : _T_11689; // @[Mux.scala 46:16:@10151.4]
  assign _T_11692 = 5'h1a == _T_10211_28; // @[Mux.scala 46:19:@10152.4]
  assign _T_11693 = _T_11692 ? _T_9260_25 : _T_11691; // @[Mux.scala 46:16:@10153.4]
  assign _T_11694 = 5'h19 == _T_10211_28; // @[Mux.scala 46:19:@10154.4]
  assign _T_11695 = _T_11694 ? _T_9260_24 : _T_11693; // @[Mux.scala 46:16:@10155.4]
  assign _T_11696 = 5'h18 == _T_10211_28; // @[Mux.scala 46:19:@10156.4]
  assign _T_11697 = _T_11696 ? _T_9260_23 : _T_11695; // @[Mux.scala 46:16:@10157.4]
  assign _T_11698 = 5'h17 == _T_10211_28; // @[Mux.scala 46:19:@10158.4]
  assign _T_11699 = _T_11698 ? _T_9260_22 : _T_11697; // @[Mux.scala 46:16:@10159.4]
  assign _T_11700 = 5'h16 == _T_10211_28; // @[Mux.scala 46:19:@10160.4]
  assign _T_11701 = _T_11700 ? _T_9260_21 : _T_11699; // @[Mux.scala 46:16:@10161.4]
  assign _T_11702 = 5'h15 == _T_10211_28; // @[Mux.scala 46:19:@10162.4]
  assign _T_11703 = _T_11702 ? _T_9260_20 : _T_11701; // @[Mux.scala 46:16:@10163.4]
  assign _T_11704 = 5'h14 == _T_10211_28; // @[Mux.scala 46:19:@10164.4]
  assign _T_11705 = _T_11704 ? _T_9260_19 : _T_11703; // @[Mux.scala 46:16:@10165.4]
  assign _T_11706 = 5'h13 == _T_10211_28; // @[Mux.scala 46:19:@10166.4]
  assign _T_11707 = _T_11706 ? _T_9260_18 : _T_11705; // @[Mux.scala 46:16:@10167.4]
  assign _T_11708 = 5'h12 == _T_10211_28; // @[Mux.scala 46:19:@10168.4]
  assign _T_11709 = _T_11708 ? _T_9260_17 : _T_11707; // @[Mux.scala 46:16:@10169.4]
  assign _T_11710 = 5'h11 == _T_10211_28; // @[Mux.scala 46:19:@10170.4]
  assign _T_11711 = _T_11710 ? _T_9260_16 : _T_11709; // @[Mux.scala 46:16:@10171.4]
  assign _T_11712 = 5'h10 == _T_10211_28; // @[Mux.scala 46:19:@10172.4]
  assign _T_11713 = _T_11712 ? _T_9260_15 : _T_11711; // @[Mux.scala 46:16:@10173.4]
  assign _T_11714 = 5'hf == _T_10211_28; // @[Mux.scala 46:19:@10174.4]
  assign _T_11715 = _T_11714 ? _T_9260_14 : _T_11713; // @[Mux.scala 46:16:@10175.4]
  assign _T_11716 = 5'he == _T_10211_28; // @[Mux.scala 46:19:@10176.4]
  assign _T_11717 = _T_11716 ? _T_9260_13 : _T_11715; // @[Mux.scala 46:16:@10177.4]
  assign _T_11718 = 5'hd == _T_10211_28; // @[Mux.scala 46:19:@10178.4]
  assign _T_11719 = _T_11718 ? _T_9260_12 : _T_11717; // @[Mux.scala 46:16:@10179.4]
  assign _T_11720 = 5'hc == _T_10211_28; // @[Mux.scala 46:19:@10180.4]
  assign _T_11721 = _T_11720 ? _T_9260_11 : _T_11719; // @[Mux.scala 46:16:@10181.4]
  assign _T_11722 = 5'hb == _T_10211_28; // @[Mux.scala 46:19:@10182.4]
  assign _T_11723 = _T_11722 ? _T_9260_10 : _T_11721; // @[Mux.scala 46:16:@10183.4]
  assign _T_11724 = 5'ha == _T_10211_28; // @[Mux.scala 46:19:@10184.4]
  assign _T_11725 = _T_11724 ? _T_9260_9 : _T_11723; // @[Mux.scala 46:16:@10185.4]
  assign _T_11726 = 5'h9 == _T_10211_28; // @[Mux.scala 46:19:@10186.4]
  assign _T_11727 = _T_11726 ? _T_9260_8 : _T_11725; // @[Mux.scala 46:16:@10187.4]
  assign _T_11728 = 5'h8 == _T_10211_28; // @[Mux.scala 46:19:@10188.4]
  assign _T_11729 = _T_11728 ? _T_9260_7 : _T_11727; // @[Mux.scala 46:16:@10189.4]
  assign _T_11730 = 5'h7 == _T_10211_28; // @[Mux.scala 46:19:@10190.4]
  assign _T_11731 = _T_11730 ? _T_9260_6 : _T_11729; // @[Mux.scala 46:16:@10191.4]
  assign _T_11732 = 5'h6 == _T_10211_28; // @[Mux.scala 46:19:@10192.4]
  assign _T_11733 = _T_11732 ? _T_9260_5 : _T_11731; // @[Mux.scala 46:16:@10193.4]
  assign _T_11734 = 5'h5 == _T_10211_28; // @[Mux.scala 46:19:@10194.4]
  assign _T_11735 = _T_11734 ? _T_9260_4 : _T_11733; // @[Mux.scala 46:16:@10195.4]
  assign _T_11736 = 5'h4 == _T_10211_28; // @[Mux.scala 46:19:@10196.4]
  assign _T_11737 = _T_11736 ? _T_9260_3 : _T_11735; // @[Mux.scala 46:16:@10197.4]
  assign _T_11738 = 5'h3 == _T_10211_28; // @[Mux.scala 46:19:@10198.4]
  assign _T_11739 = _T_11738 ? _T_9260_2 : _T_11737; // @[Mux.scala 46:16:@10199.4]
  assign _T_11740 = 5'h2 == _T_10211_28; // @[Mux.scala 46:19:@10200.4]
  assign _T_11741 = _T_11740 ? _T_9260_1 : _T_11739; // @[Mux.scala 46:16:@10201.4]
  assign _T_11742 = 5'h1 == _T_10211_28; // @[Mux.scala 46:19:@10202.4]
  assign _T_11743 = _T_11742 ? _T_9260_0 : _T_11741; // @[Mux.scala 46:16:@10203.4]
  assign _T_11775 = 5'h1e == _T_10211_29; // @[Mux.scala 46:19:@10205.4]
  assign _T_11776 = _T_11775 ? _T_9260_29 : 8'h0; // @[Mux.scala 46:16:@10206.4]
  assign _T_11777 = 5'h1d == _T_10211_29; // @[Mux.scala 46:19:@10207.4]
  assign _T_11778 = _T_11777 ? _T_9260_28 : _T_11776; // @[Mux.scala 46:16:@10208.4]
  assign _T_11779 = 5'h1c == _T_10211_29; // @[Mux.scala 46:19:@10209.4]
  assign _T_11780 = _T_11779 ? _T_9260_27 : _T_11778; // @[Mux.scala 46:16:@10210.4]
  assign _T_11781 = 5'h1b == _T_10211_29; // @[Mux.scala 46:19:@10211.4]
  assign _T_11782 = _T_11781 ? _T_9260_26 : _T_11780; // @[Mux.scala 46:16:@10212.4]
  assign _T_11783 = 5'h1a == _T_10211_29; // @[Mux.scala 46:19:@10213.4]
  assign _T_11784 = _T_11783 ? _T_9260_25 : _T_11782; // @[Mux.scala 46:16:@10214.4]
  assign _T_11785 = 5'h19 == _T_10211_29; // @[Mux.scala 46:19:@10215.4]
  assign _T_11786 = _T_11785 ? _T_9260_24 : _T_11784; // @[Mux.scala 46:16:@10216.4]
  assign _T_11787 = 5'h18 == _T_10211_29; // @[Mux.scala 46:19:@10217.4]
  assign _T_11788 = _T_11787 ? _T_9260_23 : _T_11786; // @[Mux.scala 46:16:@10218.4]
  assign _T_11789 = 5'h17 == _T_10211_29; // @[Mux.scala 46:19:@10219.4]
  assign _T_11790 = _T_11789 ? _T_9260_22 : _T_11788; // @[Mux.scala 46:16:@10220.4]
  assign _T_11791 = 5'h16 == _T_10211_29; // @[Mux.scala 46:19:@10221.4]
  assign _T_11792 = _T_11791 ? _T_9260_21 : _T_11790; // @[Mux.scala 46:16:@10222.4]
  assign _T_11793 = 5'h15 == _T_10211_29; // @[Mux.scala 46:19:@10223.4]
  assign _T_11794 = _T_11793 ? _T_9260_20 : _T_11792; // @[Mux.scala 46:16:@10224.4]
  assign _T_11795 = 5'h14 == _T_10211_29; // @[Mux.scala 46:19:@10225.4]
  assign _T_11796 = _T_11795 ? _T_9260_19 : _T_11794; // @[Mux.scala 46:16:@10226.4]
  assign _T_11797 = 5'h13 == _T_10211_29; // @[Mux.scala 46:19:@10227.4]
  assign _T_11798 = _T_11797 ? _T_9260_18 : _T_11796; // @[Mux.scala 46:16:@10228.4]
  assign _T_11799 = 5'h12 == _T_10211_29; // @[Mux.scala 46:19:@10229.4]
  assign _T_11800 = _T_11799 ? _T_9260_17 : _T_11798; // @[Mux.scala 46:16:@10230.4]
  assign _T_11801 = 5'h11 == _T_10211_29; // @[Mux.scala 46:19:@10231.4]
  assign _T_11802 = _T_11801 ? _T_9260_16 : _T_11800; // @[Mux.scala 46:16:@10232.4]
  assign _T_11803 = 5'h10 == _T_10211_29; // @[Mux.scala 46:19:@10233.4]
  assign _T_11804 = _T_11803 ? _T_9260_15 : _T_11802; // @[Mux.scala 46:16:@10234.4]
  assign _T_11805 = 5'hf == _T_10211_29; // @[Mux.scala 46:19:@10235.4]
  assign _T_11806 = _T_11805 ? _T_9260_14 : _T_11804; // @[Mux.scala 46:16:@10236.4]
  assign _T_11807 = 5'he == _T_10211_29; // @[Mux.scala 46:19:@10237.4]
  assign _T_11808 = _T_11807 ? _T_9260_13 : _T_11806; // @[Mux.scala 46:16:@10238.4]
  assign _T_11809 = 5'hd == _T_10211_29; // @[Mux.scala 46:19:@10239.4]
  assign _T_11810 = _T_11809 ? _T_9260_12 : _T_11808; // @[Mux.scala 46:16:@10240.4]
  assign _T_11811 = 5'hc == _T_10211_29; // @[Mux.scala 46:19:@10241.4]
  assign _T_11812 = _T_11811 ? _T_9260_11 : _T_11810; // @[Mux.scala 46:16:@10242.4]
  assign _T_11813 = 5'hb == _T_10211_29; // @[Mux.scala 46:19:@10243.4]
  assign _T_11814 = _T_11813 ? _T_9260_10 : _T_11812; // @[Mux.scala 46:16:@10244.4]
  assign _T_11815 = 5'ha == _T_10211_29; // @[Mux.scala 46:19:@10245.4]
  assign _T_11816 = _T_11815 ? _T_9260_9 : _T_11814; // @[Mux.scala 46:16:@10246.4]
  assign _T_11817 = 5'h9 == _T_10211_29; // @[Mux.scala 46:19:@10247.4]
  assign _T_11818 = _T_11817 ? _T_9260_8 : _T_11816; // @[Mux.scala 46:16:@10248.4]
  assign _T_11819 = 5'h8 == _T_10211_29; // @[Mux.scala 46:19:@10249.4]
  assign _T_11820 = _T_11819 ? _T_9260_7 : _T_11818; // @[Mux.scala 46:16:@10250.4]
  assign _T_11821 = 5'h7 == _T_10211_29; // @[Mux.scala 46:19:@10251.4]
  assign _T_11822 = _T_11821 ? _T_9260_6 : _T_11820; // @[Mux.scala 46:16:@10252.4]
  assign _T_11823 = 5'h6 == _T_10211_29; // @[Mux.scala 46:19:@10253.4]
  assign _T_11824 = _T_11823 ? _T_9260_5 : _T_11822; // @[Mux.scala 46:16:@10254.4]
  assign _T_11825 = 5'h5 == _T_10211_29; // @[Mux.scala 46:19:@10255.4]
  assign _T_11826 = _T_11825 ? _T_9260_4 : _T_11824; // @[Mux.scala 46:16:@10256.4]
  assign _T_11827 = 5'h4 == _T_10211_29; // @[Mux.scala 46:19:@10257.4]
  assign _T_11828 = _T_11827 ? _T_9260_3 : _T_11826; // @[Mux.scala 46:16:@10258.4]
  assign _T_11829 = 5'h3 == _T_10211_29; // @[Mux.scala 46:19:@10259.4]
  assign _T_11830 = _T_11829 ? _T_9260_2 : _T_11828; // @[Mux.scala 46:16:@10260.4]
  assign _T_11831 = 5'h2 == _T_10211_29; // @[Mux.scala 46:19:@10261.4]
  assign _T_11832 = _T_11831 ? _T_9260_1 : _T_11830; // @[Mux.scala 46:16:@10262.4]
  assign _T_11833 = 5'h1 == _T_10211_29; // @[Mux.scala 46:19:@10263.4]
  assign _T_11834 = _T_11833 ? _T_9260_0 : _T_11832; // @[Mux.scala 46:16:@10264.4]
  assign _T_11867 = 5'h1f == _T_10211_30; // @[Mux.scala 46:19:@10266.4]
  assign _T_11868 = _T_11867 ? _T_9260_30 : 8'h0; // @[Mux.scala 46:16:@10267.4]
  assign _T_11869 = 5'h1e == _T_10211_30; // @[Mux.scala 46:19:@10268.4]
  assign _T_11870 = _T_11869 ? _T_9260_29 : _T_11868; // @[Mux.scala 46:16:@10269.4]
  assign _T_11871 = 5'h1d == _T_10211_30; // @[Mux.scala 46:19:@10270.4]
  assign _T_11872 = _T_11871 ? _T_9260_28 : _T_11870; // @[Mux.scala 46:16:@10271.4]
  assign _T_11873 = 5'h1c == _T_10211_30; // @[Mux.scala 46:19:@10272.4]
  assign _T_11874 = _T_11873 ? _T_9260_27 : _T_11872; // @[Mux.scala 46:16:@10273.4]
  assign _T_11875 = 5'h1b == _T_10211_30; // @[Mux.scala 46:19:@10274.4]
  assign _T_11876 = _T_11875 ? _T_9260_26 : _T_11874; // @[Mux.scala 46:16:@10275.4]
  assign _T_11877 = 5'h1a == _T_10211_30; // @[Mux.scala 46:19:@10276.4]
  assign _T_11878 = _T_11877 ? _T_9260_25 : _T_11876; // @[Mux.scala 46:16:@10277.4]
  assign _T_11879 = 5'h19 == _T_10211_30; // @[Mux.scala 46:19:@10278.4]
  assign _T_11880 = _T_11879 ? _T_9260_24 : _T_11878; // @[Mux.scala 46:16:@10279.4]
  assign _T_11881 = 5'h18 == _T_10211_30; // @[Mux.scala 46:19:@10280.4]
  assign _T_11882 = _T_11881 ? _T_9260_23 : _T_11880; // @[Mux.scala 46:16:@10281.4]
  assign _T_11883 = 5'h17 == _T_10211_30; // @[Mux.scala 46:19:@10282.4]
  assign _T_11884 = _T_11883 ? _T_9260_22 : _T_11882; // @[Mux.scala 46:16:@10283.4]
  assign _T_11885 = 5'h16 == _T_10211_30; // @[Mux.scala 46:19:@10284.4]
  assign _T_11886 = _T_11885 ? _T_9260_21 : _T_11884; // @[Mux.scala 46:16:@10285.4]
  assign _T_11887 = 5'h15 == _T_10211_30; // @[Mux.scala 46:19:@10286.4]
  assign _T_11888 = _T_11887 ? _T_9260_20 : _T_11886; // @[Mux.scala 46:16:@10287.4]
  assign _T_11889 = 5'h14 == _T_10211_30; // @[Mux.scala 46:19:@10288.4]
  assign _T_11890 = _T_11889 ? _T_9260_19 : _T_11888; // @[Mux.scala 46:16:@10289.4]
  assign _T_11891 = 5'h13 == _T_10211_30; // @[Mux.scala 46:19:@10290.4]
  assign _T_11892 = _T_11891 ? _T_9260_18 : _T_11890; // @[Mux.scala 46:16:@10291.4]
  assign _T_11893 = 5'h12 == _T_10211_30; // @[Mux.scala 46:19:@10292.4]
  assign _T_11894 = _T_11893 ? _T_9260_17 : _T_11892; // @[Mux.scala 46:16:@10293.4]
  assign _T_11895 = 5'h11 == _T_10211_30; // @[Mux.scala 46:19:@10294.4]
  assign _T_11896 = _T_11895 ? _T_9260_16 : _T_11894; // @[Mux.scala 46:16:@10295.4]
  assign _T_11897 = 5'h10 == _T_10211_30; // @[Mux.scala 46:19:@10296.4]
  assign _T_11898 = _T_11897 ? _T_9260_15 : _T_11896; // @[Mux.scala 46:16:@10297.4]
  assign _T_11899 = 5'hf == _T_10211_30; // @[Mux.scala 46:19:@10298.4]
  assign _T_11900 = _T_11899 ? _T_9260_14 : _T_11898; // @[Mux.scala 46:16:@10299.4]
  assign _T_11901 = 5'he == _T_10211_30; // @[Mux.scala 46:19:@10300.4]
  assign _T_11902 = _T_11901 ? _T_9260_13 : _T_11900; // @[Mux.scala 46:16:@10301.4]
  assign _T_11903 = 5'hd == _T_10211_30; // @[Mux.scala 46:19:@10302.4]
  assign _T_11904 = _T_11903 ? _T_9260_12 : _T_11902; // @[Mux.scala 46:16:@10303.4]
  assign _T_11905 = 5'hc == _T_10211_30; // @[Mux.scala 46:19:@10304.4]
  assign _T_11906 = _T_11905 ? _T_9260_11 : _T_11904; // @[Mux.scala 46:16:@10305.4]
  assign _T_11907 = 5'hb == _T_10211_30; // @[Mux.scala 46:19:@10306.4]
  assign _T_11908 = _T_11907 ? _T_9260_10 : _T_11906; // @[Mux.scala 46:16:@10307.4]
  assign _T_11909 = 5'ha == _T_10211_30; // @[Mux.scala 46:19:@10308.4]
  assign _T_11910 = _T_11909 ? _T_9260_9 : _T_11908; // @[Mux.scala 46:16:@10309.4]
  assign _T_11911 = 5'h9 == _T_10211_30; // @[Mux.scala 46:19:@10310.4]
  assign _T_11912 = _T_11911 ? _T_9260_8 : _T_11910; // @[Mux.scala 46:16:@10311.4]
  assign _T_11913 = 5'h8 == _T_10211_30; // @[Mux.scala 46:19:@10312.4]
  assign _T_11914 = _T_11913 ? _T_9260_7 : _T_11912; // @[Mux.scala 46:16:@10313.4]
  assign _T_11915 = 5'h7 == _T_10211_30; // @[Mux.scala 46:19:@10314.4]
  assign _T_11916 = _T_11915 ? _T_9260_6 : _T_11914; // @[Mux.scala 46:16:@10315.4]
  assign _T_11917 = 5'h6 == _T_10211_30; // @[Mux.scala 46:19:@10316.4]
  assign _T_11918 = _T_11917 ? _T_9260_5 : _T_11916; // @[Mux.scala 46:16:@10317.4]
  assign _T_11919 = 5'h5 == _T_10211_30; // @[Mux.scala 46:19:@10318.4]
  assign _T_11920 = _T_11919 ? _T_9260_4 : _T_11918; // @[Mux.scala 46:16:@10319.4]
  assign _T_11921 = 5'h4 == _T_10211_30; // @[Mux.scala 46:19:@10320.4]
  assign _T_11922 = _T_11921 ? _T_9260_3 : _T_11920; // @[Mux.scala 46:16:@10321.4]
  assign _T_11923 = 5'h3 == _T_10211_30; // @[Mux.scala 46:19:@10322.4]
  assign _T_11924 = _T_11923 ? _T_9260_2 : _T_11922; // @[Mux.scala 46:16:@10323.4]
  assign _T_11925 = 5'h2 == _T_10211_30; // @[Mux.scala 46:19:@10324.4]
  assign _T_11926 = _T_11925 ? _T_9260_1 : _T_11924; // @[Mux.scala 46:16:@10325.4]
  assign _T_11927 = 5'h1 == _T_10211_30; // @[Mux.scala 46:19:@10326.4]
  assign _T_11928 = _T_11927 ? _T_9260_0 : _T_11926; // @[Mux.scala 46:16:@10327.4]
  assign _T_11962 = 6'h20 == _T_10211_31; // @[Mux.scala 46:19:@10329.4]
  assign _T_11963 = _T_11962 ? _T_9260_31 : 8'h0; // @[Mux.scala 46:16:@10330.4]
  assign _T_11964 = 6'h1f == _T_10211_31; // @[Mux.scala 46:19:@10331.4]
  assign _T_11965 = _T_11964 ? _T_9260_30 : _T_11963; // @[Mux.scala 46:16:@10332.4]
  assign _T_11966 = 6'h1e == _T_10211_31; // @[Mux.scala 46:19:@10333.4]
  assign _T_11967 = _T_11966 ? _T_9260_29 : _T_11965; // @[Mux.scala 46:16:@10334.4]
  assign _T_11968 = 6'h1d == _T_10211_31; // @[Mux.scala 46:19:@10335.4]
  assign _T_11969 = _T_11968 ? _T_9260_28 : _T_11967; // @[Mux.scala 46:16:@10336.4]
  assign _T_11970 = 6'h1c == _T_10211_31; // @[Mux.scala 46:19:@10337.4]
  assign _T_11971 = _T_11970 ? _T_9260_27 : _T_11969; // @[Mux.scala 46:16:@10338.4]
  assign _T_11972 = 6'h1b == _T_10211_31; // @[Mux.scala 46:19:@10339.4]
  assign _T_11973 = _T_11972 ? _T_9260_26 : _T_11971; // @[Mux.scala 46:16:@10340.4]
  assign _T_11974 = 6'h1a == _T_10211_31; // @[Mux.scala 46:19:@10341.4]
  assign _T_11975 = _T_11974 ? _T_9260_25 : _T_11973; // @[Mux.scala 46:16:@10342.4]
  assign _T_11976 = 6'h19 == _T_10211_31; // @[Mux.scala 46:19:@10343.4]
  assign _T_11977 = _T_11976 ? _T_9260_24 : _T_11975; // @[Mux.scala 46:16:@10344.4]
  assign _T_11978 = 6'h18 == _T_10211_31; // @[Mux.scala 46:19:@10345.4]
  assign _T_11979 = _T_11978 ? _T_9260_23 : _T_11977; // @[Mux.scala 46:16:@10346.4]
  assign _T_11980 = 6'h17 == _T_10211_31; // @[Mux.scala 46:19:@10347.4]
  assign _T_11981 = _T_11980 ? _T_9260_22 : _T_11979; // @[Mux.scala 46:16:@10348.4]
  assign _T_11982 = 6'h16 == _T_10211_31; // @[Mux.scala 46:19:@10349.4]
  assign _T_11983 = _T_11982 ? _T_9260_21 : _T_11981; // @[Mux.scala 46:16:@10350.4]
  assign _T_11984 = 6'h15 == _T_10211_31; // @[Mux.scala 46:19:@10351.4]
  assign _T_11985 = _T_11984 ? _T_9260_20 : _T_11983; // @[Mux.scala 46:16:@10352.4]
  assign _T_11986 = 6'h14 == _T_10211_31; // @[Mux.scala 46:19:@10353.4]
  assign _T_11987 = _T_11986 ? _T_9260_19 : _T_11985; // @[Mux.scala 46:16:@10354.4]
  assign _T_11988 = 6'h13 == _T_10211_31; // @[Mux.scala 46:19:@10355.4]
  assign _T_11989 = _T_11988 ? _T_9260_18 : _T_11987; // @[Mux.scala 46:16:@10356.4]
  assign _T_11990 = 6'h12 == _T_10211_31; // @[Mux.scala 46:19:@10357.4]
  assign _T_11991 = _T_11990 ? _T_9260_17 : _T_11989; // @[Mux.scala 46:16:@10358.4]
  assign _T_11992 = 6'h11 == _T_10211_31; // @[Mux.scala 46:19:@10359.4]
  assign _T_11993 = _T_11992 ? _T_9260_16 : _T_11991; // @[Mux.scala 46:16:@10360.4]
  assign _T_11994 = 6'h10 == _T_10211_31; // @[Mux.scala 46:19:@10361.4]
  assign _T_11995 = _T_11994 ? _T_9260_15 : _T_11993; // @[Mux.scala 46:16:@10362.4]
  assign _T_11996 = 6'hf == _T_10211_31; // @[Mux.scala 46:19:@10363.4]
  assign _T_11997 = _T_11996 ? _T_9260_14 : _T_11995; // @[Mux.scala 46:16:@10364.4]
  assign _T_11998 = 6'he == _T_10211_31; // @[Mux.scala 46:19:@10365.4]
  assign _T_11999 = _T_11998 ? _T_9260_13 : _T_11997; // @[Mux.scala 46:16:@10366.4]
  assign _T_12000 = 6'hd == _T_10211_31; // @[Mux.scala 46:19:@10367.4]
  assign _T_12001 = _T_12000 ? _T_9260_12 : _T_11999; // @[Mux.scala 46:16:@10368.4]
  assign _T_12002 = 6'hc == _T_10211_31; // @[Mux.scala 46:19:@10369.4]
  assign _T_12003 = _T_12002 ? _T_9260_11 : _T_12001; // @[Mux.scala 46:16:@10370.4]
  assign _T_12004 = 6'hb == _T_10211_31; // @[Mux.scala 46:19:@10371.4]
  assign _T_12005 = _T_12004 ? _T_9260_10 : _T_12003; // @[Mux.scala 46:16:@10372.4]
  assign _T_12006 = 6'ha == _T_10211_31; // @[Mux.scala 46:19:@10373.4]
  assign _T_12007 = _T_12006 ? _T_9260_9 : _T_12005; // @[Mux.scala 46:16:@10374.4]
  assign _T_12008 = 6'h9 == _T_10211_31; // @[Mux.scala 46:19:@10375.4]
  assign _T_12009 = _T_12008 ? _T_9260_8 : _T_12007; // @[Mux.scala 46:16:@10376.4]
  assign _T_12010 = 6'h8 == _T_10211_31; // @[Mux.scala 46:19:@10377.4]
  assign _T_12011 = _T_12010 ? _T_9260_7 : _T_12009; // @[Mux.scala 46:16:@10378.4]
  assign _T_12012 = 6'h7 == _T_10211_31; // @[Mux.scala 46:19:@10379.4]
  assign _T_12013 = _T_12012 ? _T_9260_6 : _T_12011; // @[Mux.scala 46:16:@10380.4]
  assign _T_12014 = 6'h6 == _T_10211_31; // @[Mux.scala 46:19:@10381.4]
  assign _T_12015 = _T_12014 ? _T_9260_5 : _T_12013; // @[Mux.scala 46:16:@10382.4]
  assign _T_12016 = 6'h5 == _T_10211_31; // @[Mux.scala 46:19:@10383.4]
  assign _T_12017 = _T_12016 ? _T_9260_4 : _T_12015; // @[Mux.scala 46:16:@10384.4]
  assign _T_12018 = 6'h4 == _T_10211_31; // @[Mux.scala 46:19:@10385.4]
  assign _T_12019 = _T_12018 ? _T_9260_3 : _T_12017; // @[Mux.scala 46:16:@10386.4]
  assign _T_12020 = 6'h3 == _T_10211_31; // @[Mux.scala 46:19:@10387.4]
  assign _T_12021 = _T_12020 ? _T_9260_2 : _T_12019; // @[Mux.scala 46:16:@10388.4]
  assign _T_12022 = 6'h2 == _T_10211_31; // @[Mux.scala 46:19:@10389.4]
  assign _T_12023 = _T_12022 ? _T_9260_1 : _T_12021; // @[Mux.scala 46:16:@10390.4]
  assign _T_12024 = 6'h1 == _T_10211_31; // @[Mux.scala 46:19:@10391.4]
  assign _T_12025 = _T_12024 ? _T_9260_0 : _T_12023; // @[Mux.scala 46:16:@10392.4]
  assign _T_12060 = 6'h21 == _T_10211_32; // @[Mux.scala 46:19:@10394.4]
  assign _T_12061 = _T_12060 ? _T_9260_32 : 8'h0; // @[Mux.scala 46:16:@10395.4]
  assign _T_12062 = 6'h20 == _T_10211_32; // @[Mux.scala 46:19:@10396.4]
  assign _T_12063 = _T_12062 ? _T_9260_31 : _T_12061; // @[Mux.scala 46:16:@10397.4]
  assign _T_12064 = 6'h1f == _T_10211_32; // @[Mux.scala 46:19:@10398.4]
  assign _T_12065 = _T_12064 ? _T_9260_30 : _T_12063; // @[Mux.scala 46:16:@10399.4]
  assign _T_12066 = 6'h1e == _T_10211_32; // @[Mux.scala 46:19:@10400.4]
  assign _T_12067 = _T_12066 ? _T_9260_29 : _T_12065; // @[Mux.scala 46:16:@10401.4]
  assign _T_12068 = 6'h1d == _T_10211_32; // @[Mux.scala 46:19:@10402.4]
  assign _T_12069 = _T_12068 ? _T_9260_28 : _T_12067; // @[Mux.scala 46:16:@10403.4]
  assign _T_12070 = 6'h1c == _T_10211_32; // @[Mux.scala 46:19:@10404.4]
  assign _T_12071 = _T_12070 ? _T_9260_27 : _T_12069; // @[Mux.scala 46:16:@10405.4]
  assign _T_12072 = 6'h1b == _T_10211_32; // @[Mux.scala 46:19:@10406.4]
  assign _T_12073 = _T_12072 ? _T_9260_26 : _T_12071; // @[Mux.scala 46:16:@10407.4]
  assign _T_12074 = 6'h1a == _T_10211_32; // @[Mux.scala 46:19:@10408.4]
  assign _T_12075 = _T_12074 ? _T_9260_25 : _T_12073; // @[Mux.scala 46:16:@10409.4]
  assign _T_12076 = 6'h19 == _T_10211_32; // @[Mux.scala 46:19:@10410.4]
  assign _T_12077 = _T_12076 ? _T_9260_24 : _T_12075; // @[Mux.scala 46:16:@10411.4]
  assign _T_12078 = 6'h18 == _T_10211_32; // @[Mux.scala 46:19:@10412.4]
  assign _T_12079 = _T_12078 ? _T_9260_23 : _T_12077; // @[Mux.scala 46:16:@10413.4]
  assign _T_12080 = 6'h17 == _T_10211_32; // @[Mux.scala 46:19:@10414.4]
  assign _T_12081 = _T_12080 ? _T_9260_22 : _T_12079; // @[Mux.scala 46:16:@10415.4]
  assign _T_12082 = 6'h16 == _T_10211_32; // @[Mux.scala 46:19:@10416.4]
  assign _T_12083 = _T_12082 ? _T_9260_21 : _T_12081; // @[Mux.scala 46:16:@10417.4]
  assign _T_12084 = 6'h15 == _T_10211_32; // @[Mux.scala 46:19:@10418.4]
  assign _T_12085 = _T_12084 ? _T_9260_20 : _T_12083; // @[Mux.scala 46:16:@10419.4]
  assign _T_12086 = 6'h14 == _T_10211_32; // @[Mux.scala 46:19:@10420.4]
  assign _T_12087 = _T_12086 ? _T_9260_19 : _T_12085; // @[Mux.scala 46:16:@10421.4]
  assign _T_12088 = 6'h13 == _T_10211_32; // @[Mux.scala 46:19:@10422.4]
  assign _T_12089 = _T_12088 ? _T_9260_18 : _T_12087; // @[Mux.scala 46:16:@10423.4]
  assign _T_12090 = 6'h12 == _T_10211_32; // @[Mux.scala 46:19:@10424.4]
  assign _T_12091 = _T_12090 ? _T_9260_17 : _T_12089; // @[Mux.scala 46:16:@10425.4]
  assign _T_12092 = 6'h11 == _T_10211_32; // @[Mux.scala 46:19:@10426.4]
  assign _T_12093 = _T_12092 ? _T_9260_16 : _T_12091; // @[Mux.scala 46:16:@10427.4]
  assign _T_12094 = 6'h10 == _T_10211_32; // @[Mux.scala 46:19:@10428.4]
  assign _T_12095 = _T_12094 ? _T_9260_15 : _T_12093; // @[Mux.scala 46:16:@10429.4]
  assign _T_12096 = 6'hf == _T_10211_32; // @[Mux.scala 46:19:@10430.4]
  assign _T_12097 = _T_12096 ? _T_9260_14 : _T_12095; // @[Mux.scala 46:16:@10431.4]
  assign _T_12098 = 6'he == _T_10211_32; // @[Mux.scala 46:19:@10432.4]
  assign _T_12099 = _T_12098 ? _T_9260_13 : _T_12097; // @[Mux.scala 46:16:@10433.4]
  assign _T_12100 = 6'hd == _T_10211_32; // @[Mux.scala 46:19:@10434.4]
  assign _T_12101 = _T_12100 ? _T_9260_12 : _T_12099; // @[Mux.scala 46:16:@10435.4]
  assign _T_12102 = 6'hc == _T_10211_32; // @[Mux.scala 46:19:@10436.4]
  assign _T_12103 = _T_12102 ? _T_9260_11 : _T_12101; // @[Mux.scala 46:16:@10437.4]
  assign _T_12104 = 6'hb == _T_10211_32; // @[Mux.scala 46:19:@10438.4]
  assign _T_12105 = _T_12104 ? _T_9260_10 : _T_12103; // @[Mux.scala 46:16:@10439.4]
  assign _T_12106 = 6'ha == _T_10211_32; // @[Mux.scala 46:19:@10440.4]
  assign _T_12107 = _T_12106 ? _T_9260_9 : _T_12105; // @[Mux.scala 46:16:@10441.4]
  assign _T_12108 = 6'h9 == _T_10211_32; // @[Mux.scala 46:19:@10442.4]
  assign _T_12109 = _T_12108 ? _T_9260_8 : _T_12107; // @[Mux.scala 46:16:@10443.4]
  assign _T_12110 = 6'h8 == _T_10211_32; // @[Mux.scala 46:19:@10444.4]
  assign _T_12111 = _T_12110 ? _T_9260_7 : _T_12109; // @[Mux.scala 46:16:@10445.4]
  assign _T_12112 = 6'h7 == _T_10211_32; // @[Mux.scala 46:19:@10446.4]
  assign _T_12113 = _T_12112 ? _T_9260_6 : _T_12111; // @[Mux.scala 46:16:@10447.4]
  assign _T_12114 = 6'h6 == _T_10211_32; // @[Mux.scala 46:19:@10448.4]
  assign _T_12115 = _T_12114 ? _T_9260_5 : _T_12113; // @[Mux.scala 46:16:@10449.4]
  assign _T_12116 = 6'h5 == _T_10211_32; // @[Mux.scala 46:19:@10450.4]
  assign _T_12117 = _T_12116 ? _T_9260_4 : _T_12115; // @[Mux.scala 46:16:@10451.4]
  assign _T_12118 = 6'h4 == _T_10211_32; // @[Mux.scala 46:19:@10452.4]
  assign _T_12119 = _T_12118 ? _T_9260_3 : _T_12117; // @[Mux.scala 46:16:@10453.4]
  assign _T_12120 = 6'h3 == _T_10211_32; // @[Mux.scala 46:19:@10454.4]
  assign _T_12121 = _T_12120 ? _T_9260_2 : _T_12119; // @[Mux.scala 46:16:@10455.4]
  assign _T_12122 = 6'h2 == _T_10211_32; // @[Mux.scala 46:19:@10456.4]
  assign _T_12123 = _T_12122 ? _T_9260_1 : _T_12121; // @[Mux.scala 46:16:@10457.4]
  assign _T_12124 = 6'h1 == _T_10211_32; // @[Mux.scala 46:19:@10458.4]
  assign _T_12125 = _T_12124 ? _T_9260_0 : _T_12123; // @[Mux.scala 46:16:@10459.4]
  assign _T_12161 = 6'h22 == _T_10211_33; // @[Mux.scala 46:19:@10461.4]
  assign _T_12162 = _T_12161 ? _T_9260_33 : 8'h0; // @[Mux.scala 46:16:@10462.4]
  assign _T_12163 = 6'h21 == _T_10211_33; // @[Mux.scala 46:19:@10463.4]
  assign _T_12164 = _T_12163 ? _T_9260_32 : _T_12162; // @[Mux.scala 46:16:@10464.4]
  assign _T_12165 = 6'h20 == _T_10211_33; // @[Mux.scala 46:19:@10465.4]
  assign _T_12166 = _T_12165 ? _T_9260_31 : _T_12164; // @[Mux.scala 46:16:@10466.4]
  assign _T_12167 = 6'h1f == _T_10211_33; // @[Mux.scala 46:19:@10467.4]
  assign _T_12168 = _T_12167 ? _T_9260_30 : _T_12166; // @[Mux.scala 46:16:@10468.4]
  assign _T_12169 = 6'h1e == _T_10211_33; // @[Mux.scala 46:19:@10469.4]
  assign _T_12170 = _T_12169 ? _T_9260_29 : _T_12168; // @[Mux.scala 46:16:@10470.4]
  assign _T_12171 = 6'h1d == _T_10211_33; // @[Mux.scala 46:19:@10471.4]
  assign _T_12172 = _T_12171 ? _T_9260_28 : _T_12170; // @[Mux.scala 46:16:@10472.4]
  assign _T_12173 = 6'h1c == _T_10211_33; // @[Mux.scala 46:19:@10473.4]
  assign _T_12174 = _T_12173 ? _T_9260_27 : _T_12172; // @[Mux.scala 46:16:@10474.4]
  assign _T_12175 = 6'h1b == _T_10211_33; // @[Mux.scala 46:19:@10475.4]
  assign _T_12176 = _T_12175 ? _T_9260_26 : _T_12174; // @[Mux.scala 46:16:@10476.4]
  assign _T_12177 = 6'h1a == _T_10211_33; // @[Mux.scala 46:19:@10477.4]
  assign _T_12178 = _T_12177 ? _T_9260_25 : _T_12176; // @[Mux.scala 46:16:@10478.4]
  assign _T_12179 = 6'h19 == _T_10211_33; // @[Mux.scala 46:19:@10479.4]
  assign _T_12180 = _T_12179 ? _T_9260_24 : _T_12178; // @[Mux.scala 46:16:@10480.4]
  assign _T_12181 = 6'h18 == _T_10211_33; // @[Mux.scala 46:19:@10481.4]
  assign _T_12182 = _T_12181 ? _T_9260_23 : _T_12180; // @[Mux.scala 46:16:@10482.4]
  assign _T_12183 = 6'h17 == _T_10211_33; // @[Mux.scala 46:19:@10483.4]
  assign _T_12184 = _T_12183 ? _T_9260_22 : _T_12182; // @[Mux.scala 46:16:@10484.4]
  assign _T_12185 = 6'h16 == _T_10211_33; // @[Mux.scala 46:19:@10485.4]
  assign _T_12186 = _T_12185 ? _T_9260_21 : _T_12184; // @[Mux.scala 46:16:@10486.4]
  assign _T_12187 = 6'h15 == _T_10211_33; // @[Mux.scala 46:19:@10487.4]
  assign _T_12188 = _T_12187 ? _T_9260_20 : _T_12186; // @[Mux.scala 46:16:@10488.4]
  assign _T_12189 = 6'h14 == _T_10211_33; // @[Mux.scala 46:19:@10489.4]
  assign _T_12190 = _T_12189 ? _T_9260_19 : _T_12188; // @[Mux.scala 46:16:@10490.4]
  assign _T_12191 = 6'h13 == _T_10211_33; // @[Mux.scala 46:19:@10491.4]
  assign _T_12192 = _T_12191 ? _T_9260_18 : _T_12190; // @[Mux.scala 46:16:@10492.4]
  assign _T_12193 = 6'h12 == _T_10211_33; // @[Mux.scala 46:19:@10493.4]
  assign _T_12194 = _T_12193 ? _T_9260_17 : _T_12192; // @[Mux.scala 46:16:@10494.4]
  assign _T_12195 = 6'h11 == _T_10211_33; // @[Mux.scala 46:19:@10495.4]
  assign _T_12196 = _T_12195 ? _T_9260_16 : _T_12194; // @[Mux.scala 46:16:@10496.4]
  assign _T_12197 = 6'h10 == _T_10211_33; // @[Mux.scala 46:19:@10497.4]
  assign _T_12198 = _T_12197 ? _T_9260_15 : _T_12196; // @[Mux.scala 46:16:@10498.4]
  assign _T_12199 = 6'hf == _T_10211_33; // @[Mux.scala 46:19:@10499.4]
  assign _T_12200 = _T_12199 ? _T_9260_14 : _T_12198; // @[Mux.scala 46:16:@10500.4]
  assign _T_12201 = 6'he == _T_10211_33; // @[Mux.scala 46:19:@10501.4]
  assign _T_12202 = _T_12201 ? _T_9260_13 : _T_12200; // @[Mux.scala 46:16:@10502.4]
  assign _T_12203 = 6'hd == _T_10211_33; // @[Mux.scala 46:19:@10503.4]
  assign _T_12204 = _T_12203 ? _T_9260_12 : _T_12202; // @[Mux.scala 46:16:@10504.4]
  assign _T_12205 = 6'hc == _T_10211_33; // @[Mux.scala 46:19:@10505.4]
  assign _T_12206 = _T_12205 ? _T_9260_11 : _T_12204; // @[Mux.scala 46:16:@10506.4]
  assign _T_12207 = 6'hb == _T_10211_33; // @[Mux.scala 46:19:@10507.4]
  assign _T_12208 = _T_12207 ? _T_9260_10 : _T_12206; // @[Mux.scala 46:16:@10508.4]
  assign _T_12209 = 6'ha == _T_10211_33; // @[Mux.scala 46:19:@10509.4]
  assign _T_12210 = _T_12209 ? _T_9260_9 : _T_12208; // @[Mux.scala 46:16:@10510.4]
  assign _T_12211 = 6'h9 == _T_10211_33; // @[Mux.scala 46:19:@10511.4]
  assign _T_12212 = _T_12211 ? _T_9260_8 : _T_12210; // @[Mux.scala 46:16:@10512.4]
  assign _T_12213 = 6'h8 == _T_10211_33; // @[Mux.scala 46:19:@10513.4]
  assign _T_12214 = _T_12213 ? _T_9260_7 : _T_12212; // @[Mux.scala 46:16:@10514.4]
  assign _T_12215 = 6'h7 == _T_10211_33; // @[Mux.scala 46:19:@10515.4]
  assign _T_12216 = _T_12215 ? _T_9260_6 : _T_12214; // @[Mux.scala 46:16:@10516.4]
  assign _T_12217 = 6'h6 == _T_10211_33; // @[Mux.scala 46:19:@10517.4]
  assign _T_12218 = _T_12217 ? _T_9260_5 : _T_12216; // @[Mux.scala 46:16:@10518.4]
  assign _T_12219 = 6'h5 == _T_10211_33; // @[Mux.scala 46:19:@10519.4]
  assign _T_12220 = _T_12219 ? _T_9260_4 : _T_12218; // @[Mux.scala 46:16:@10520.4]
  assign _T_12221 = 6'h4 == _T_10211_33; // @[Mux.scala 46:19:@10521.4]
  assign _T_12222 = _T_12221 ? _T_9260_3 : _T_12220; // @[Mux.scala 46:16:@10522.4]
  assign _T_12223 = 6'h3 == _T_10211_33; // @[Mux.scala 46:19:@10523.4]
  assign _T_12224 = _T_12223 ? _T_9260_2 : _T_12222; // @[Mux.scala 46:16:@10524.4]
  assign _T_12225 = 6'h2 == _T_10211_33; // @[Mux.scala 46:19:@10525.4]
  assign _T_12226 = _T_12225 ? _T_9260_1 : _T_12224; // @[Mux.scala 46:16:@10526.4]
  assign _T_12227 = 6'h1 == _T_10211_33; // @[Mux.scala 46:19:@10527.4]
  assign _T_12228 = _T_12227 ? _T_9260_0 : _T_12226; // @[Mux.scala 46:16:@10528.4]
  assign _T_12265 = 6'h23 == _T_10211_34; // @[Mux.scala 46:19:@10530.4]
  assign _T_12266 = _T_12265 ? _T_9260_34 : 8'h0; // @[Mux.scala 46:16:@10531.4]
  assign _T_12267 = 6'h22 == _T_10211_34; // @[Mux.scala 46:19:@10532.4]
  assign _T_12268 = _T_12267 ? _T_9260_33 : _T_12266; // @[Mux.scala 46:16:@10533.4]
  assign _T_12269 = 6'h21 == _T_10211_34; // @[Mux.scala 46:19:@10534.4]
  assign _T_12270 = _T_12269 ? _T_9260_32 : _T_12268; // @[Mux.scala 46:16:@10535.4]
  assign _T_12271 = 6'h20 == _T_10211_34; // @[Mux.scala 46:19:@10536.4]
  assign _T_12272 = _T_12271 ? _T_9260_31 : _T_12270; // @[Mux.scala 46:16:@10537.4]
  assign _T_12273 = 6'h1f == _T_10211_34; // @[Mux.scala 46:19:@10538.4]
  assign _T_12274 = _T_12273 ? _T_9260_30 : _T_12272; // @[Mux.scala 46:16:@10539.4]
  assign _T_12275 = 6'h1e == _T_10211_34; // @[Mux.scala 46:19:@10540.4]
  assign _T_12276 = _T_12275 ? _T_9260_29 : _T_12274; // @[Mux.scala 46:16:@10541.4]
  assign _T_12277 = 6'h1d == _T_10211_34; // @[Mux.scala 46:19:@10542.4]
  assign _T_12278 = _T_12277 ? _T_9260_28 : _T_12276; // @[Mux.scala 46:16:@10543.4]
  assign _T_12279 = 6'h1c == _T_10211_34; // @[Mux.scala 46:19:@10544.4]
  assign _T_12280 = _T_12279 ? _T_9260_27 : _T_12278; // @[Mux.scala 46:16:@10545.4]
  assign _T_12281 = 6'h1b == _T_10211_34; // @[Mux.scala 46:19:@10546.4]
  assign _T_12282 = _T_12281 ? _T_9260_26 : _T_12280; // @[Mux.scala 46:16:@10547.4]
  assign _T_12283 = 6'h1a == _T_10211_34; // @[Mux.scala 46:19:@10548.4]
  assign _T_12284 = _T_12283 ? _T_9260_25 : _T_12282; // @[Mux.scala 46:16:@10549.4]
  assign _T_12285 = 6'h19 == _T_10211_34; // @[Mux.scala 46:19:@10550.4]
  assign _T_12286 = _T_12285 ? _T_9260_24 : _T_12284; // @[Mux.scala 46:16:@10551.4]
  assign _T_12287 = 6'h18 == _T_10211_34; // @[Mux.scala 46:19:@10552.4]
  assign _T_12288 = _T_12287 ? _T_9260_23 : _T_12286; // @[Mux.scala 46:16:@10553.4]
  assign _T_12289 = 6'h17 == _T_10211_34; // @[Mux.scala 46:19:@10554.4]
  assign _T_12290 = _T_12289 ? _T_9260_22 : _T_12288; // @[Mux.scala 46:16:@10555.4]
  assign _T_12291 = 6'h16 == _T_10211_34; // @[Mux.scala 46:19:@10556.4]
  assign _T_12292 = _T_12291 ? _T_9260_21 : _T_12290; // @[Mux.scala 46:16:@10557.4]
  assign _T_12293 = 6'h15 == _T_10211_34; // @[Mux.scala 46:19:@10558.4]
  assign _T_12294 = _T_12293 ? _T_9260_20 : _T_12292; // @[Mux.scala 46:16:@10559.4]
  assign _T_12295 = 6'h14 == _T_10211_34; // @[Mux.scala 46:19:@10560.4]
  assign _T_12296 = _T_12295 ? _T_9260_19 : _T_12294; // @[Mux.scala 46:16:@10561.4]
  assign _T_12297 = 6'h13 == _T_10211_34; // @[Mux.scala 46:19:@10562.4]
  assign _T_12298 = _T_12297 ? _T_9260_18 : _T_12296; // @[Mux.scala 46:16:@10563.4]
  assign _T_12299 = 6'h12 == _T_10211_34; // @[Mux.scala 46:19:@10564.4]
  assign _T_12300 = _T_12299 ? _T_9260_17 : _T_12298; // @[Mux.scala 46:16:@10565.4]
  assign _T_12301 = 6'h11 == _T_10211_34; // @[Mux.scala 46:19:@10566.4]
  assign _T_12302 = _T_12301 ? _T_9260_16 : _T_12300; // @[Mux.scala 46:16:@10567.4]
  assign _T_12303 = 6'h10 == _T_10211_34; // @[Mux.scala 46:19:@10568.4]
  assign _T_12304 = _T_12303 ? _T_9260_15 : _T_12302; // @[Mux.scala 46:16:@10569.4]
  assign _T_12305 = 6'hf == _T_10211_34; // @[Mux.scala 46:19:@10570.4]
  assign _T_12306 = _T_12305 ? _T_9260_14 : _T_12304; // @[Mux.scala 46:16:@10571.4]
  assign _T_12307 = 6'he == _T_10211_34; // @[Mux.scala 46:19:@10572.4]
  assign _T_12308 = _T_12307 ? _T_9260_13 : _T_12306; // @[Mux.scala 46:16:@10573.4]
  assign _T_12309 = 6'hd == _T_10211_34; // @[Mux.scala 46:19:@10574.4]
  assign _T_12310 = _T_12309 ? _T_9260_12 : _T_12308; // @[Mux.scala 46:16:@10575.4]
  assign _T_12311 = 6'hc == _T_10211_34; // @[Mux.scala 46:19:@10576.4]
  assign _T_12312 = _T_12311 ? _T_9260_11 : _T_12310; // @[Mux.scala 46:16:@10577.4]
  assign _T_12313 = 6'hb == _T_10211_34; // @[Mux.scala 46:19:@10578.4]
  assign _T_12314 = _T_12313 ? _T_9260_10 : _T_12312; // @[Mux.scala 46:16:@10579.4]
  assign _T_12315 = 6'ha == _T_10211_34; // @[Mux.scala 46:19:@10580.4]
  assign _T_12316 = _T_12315 ? _T_9260_9 : _T_12314; // @[Mux.scala 46:16:@10581.4]
  assign _T_12317 = 6'h9 == _T_10211_34; // @[Mux.scala 46:19:@10582.4]
  assign _T_12318 = _T_12317 ? _T_9260_8 : _T_12316; // @[Mux.scala 46:16:@10583.4]
  assign _T_12319 = 6'h8 == _T_10211_34; // @[Mux.scala 46:19:@10584.4]
  assign _T_12320 = _T_12319 ? _T_9260_7 : _T_12318; // @[Mux.scala 46:16:@10585.4]
  assign _T_12321 = 6'h7 == _T_10211_34; // @[Mux.scala 46:19:@10586.4]
  assign _T_12322 = _T_12321 ? _T_9260_6 : _T_12320; // @[Mux.scala 46:16:@10587.4]
  assign _T_12323 = 6'h6 == _T_10211_34; // @[Mux.scala 46:19:@10588.4]
  assign _T_12324 = _T_12323 ? _T_9260_5 : _T_12322; // @[Mux.scala 46:16:@10589.4]
  assign _T_12325 = 6'h5 == _T_10211_34; // @[Mux.scala 46:19:@10590.4]
  assign _T_12326 = _T_12325 ? _T_9260_4 : _T_12324; // @[Mux.scala 46:16:@10591.4]
  assign _T_12327 = 6'h4 == _T_10211_34; // @[Mux.scala 46:19:@10592.4]
  assign _T_12328 = _T_12327 ? _T_9260_3 : _T_12326; // @[Mux.scala 46:16:@10593.4]
  assign _T_12329 = 6'h3 == _T_10211_34; // @[Mux.scala 46:19:@10594.4]
  assign _T_12330 = _T_12329 ? _T_9260_2 : _T_12328; // @[Mux.scala 46:16:@10595.4]
  assign _T_12331 = 6'h2 == _T_10211_34; // @[Mux.scala 46:19:@10596.4]
  assign _T_12332 = _T_12331 ? _T_9260_1 : _T_12330; // @[Mux.scala 46:16:@10597.4]
  assign _T_12333 = 6'h1 == _T_10211_34; // @[Mux.scala 46:19:@10598.4]
  assign _T_12334 = _T_12333 ? _T_9260_0 : _T_12332; // @[Mux.scala 46:16:@10599.4]
  assign _T_12372 = 6'h24 == _T_10211_35; // @[Mux.scala 46:19:@10601.4]
  assign _T_12373 = _T_12372 ? _T_9260_35 : 8'h0; // @[Mux.scala 46:16:@10602.4]
  assign _T_12374 = 6'h23 == _T_10211_35; // @[Mux.scala 46:19:@10603.4]
  assign _T_12375 = _T_12374 ? _T_9260_34 : _T_12373; // @[Mux.scala 46:16:@10604.4]
  assign _T_12376 = 6'h22 == _T_10211_35; // @[Mux.scala 46:19:@10605.4]
  assign _T_12377 = _T_12376 ? _T_9260_33 : _T_12375; // @[Mux.scala 46:16:@10606.4]
  assign _T_12378 = 6'h21 == _T_10211_35; // @[Mux.scala 46:19:@10607.4]
  assign _T_12379 = _T_12378 ? _T_9260_32 : _T_12377; // @[Mux.scala 46:16:@10608.4]
  assign _T_12380 = 6'h20 == _T_10211_35; // @[Mux.scala 46:19:@10609.4]
  assign _T_12381 = _T_12380 ? _T_9260_31 : _T_12379; // @[Mux.scala 46:16:@10610.4]
  assign _T_12382 = 6'h1f == _T_10211_35; // @[Mux.scala 46:19:@10611.4]
  assign _T_12383 = _T_12382 ? _T_9260_30 : _T_12381; // @[Mux.scala 46:16:@10612.4]
  assign _T_12384 = 6'h1e == _T_10211_35; // @[Mux.scala 46:19:@10613.4]
  assign _T_12385 = _T_12384 ? _T_9260_29 : _T_12383; // @[Mux.scala 46:16:@10614.4]
  assign _T_12386 = 6'h1d == _T_10211_35; // @[Mux.scala 46:19:@10615.4]
  assign _T_12387 = _T_12386 ? _T_9260_28 : _T_12385; // @[Mux.scala 46:16:@10616.4]
  assign _T_12388 = 6'h1c == _T_10211_35; // @[Mux.scala 46:19:@10617.4]
  assign _T_12389 = _T_12388 ? _T_9260_27 : _T_12387; // @[Mux.scala 46:16:@10618.4]
  assign _T_12390 = 6'h1b == _T_10211_35; // @[Mux.scala 46:19:@10619.4]
  assign _T_12391 = _T_12390 ? _T_9260_26 : _T_12389; // @[Mux.scala 46:16:@10620.4]
  assign _T_12392 = 6'h1a == _T_10211_35; // @[Mux.scala 46:19:@10621.4]
  assign _T_12393 = _T_12392 ? _T_9260_25 : _T_12391; // @[Mux.scala 46:16:@10622.4]
  assign _T_12394 = 6'h19 == _T_10211_35; // @[Mux.scala 46:19:@10623.4]
  assign _T_12395 = _T_12394 ? _T_9260_24 : _T_12393; // @[Mux.scala 46:16:@10624.4]
  assign _T_12396 = 6'h18 == _T_10211_35; // @[Mux.scala 46:19:@10625.4]
  assign _T_12397 = _T_12396 ? _T_9260_23 : _T_12395; // @[Mux.scala 46:16:@10626.4]
  assign _T_12398 = 6'h17 == _T_10211_35; // @[Mux.scala 46:19:@10627.4]
  assign _T_12399 = _T_12398 ? _T_9260_22 : _T_12397; // @[Mux.scala 46:16:@10628.4]
  assign _T_12400 = 6'h16 == _T_10211_35; // @[Mux.scala 46:19:@10629.4]
  assign _T_12401 = _T_12400 ? _T_9260_21 : _T_12399; // @[Mux.scala 46:16:@10630.4]
  assign _T_12402 = 6'h15 == _T_10211_35; // @[Mux.scala 46:19:@10631.4]
  assign _T_12403 = _T_12402 ? _T_9260_20 : _T_12401; // @[Mux.scala 46:16:@10632.4]
  assign _T_12404 = 6'h14 == _T_10211_35; // @[Mux.scala 46:19:@10633.4]
  assign _T_12405 = _T_12404 ? _T_9260_19 : _T_12403; // @[Mux.scala 46:16:@10634.4]
  assign _T_12406 = 6'h13 == _T_10211_35; // @[Mux.scala 46:19:@10635.4]
  assign _T_12407 = _T_12406 ? _T_9260_18 : _T_12405; // @[Mux.scala 46:16:@10636.4]
  assign _T_12408 = 6'h12 == _T_10211_35; // @[Mux.scala 46:19:@10637.4]
  assign _T_12409 = _T_12408 ? _T_9260_17 : _T_12407; // @[Mux.scala 46:16:@10638.4]
  assign _T_12410 = 6'h11 == _T_10211_35; // @[Mux.scala 46:19:@10639.4]
  assign _T_12411 = _T_12410 ? _T_9260_16 : _T_12409; // @[Mux.scala 46:16:@10640.4]
  assign _T_12412 = 6'h10 == _T_10211_35; // @[Mux.scala 46:19:@10641.4]
  assign _T_12413 = _T_12412 ? _T_9260_15 : _T_12411; // @[Mux.scala 46:16:@10642.4]
  assign _T_12414 = 6'hf == _T_10211_35; // @[Mux.scala 46:19:@10643.4]
  assign _T_12415 = _T_12414 ? _T_9260_14 : _T_12413; // @[Mux.scala 46:16:@10644.4]
  assign _T_12416 = 6'he == _T_10211_35; // @[Mux.scala 46:19:@10645.4]
  assign _T_12417 = _T_12416 ? _T_9260_13 : _T_12415; // @[Mux.scala 46:16:@10646.4]
  assign _T_12418 = 6'hd == _T_10211_35; // @[Mux.scala 46:19:@10647.4]
  assign _T_12419 = _T_12418 ? _T_9260_12 : _T_12417; // @[Mux.scala 46:16:@10648.4]
  assign _T_12420 = 6'hc == _T_10211_35; // @[Mux.scala 46:19:@10649.4]
  assign _T_12421 = _T_12420 ? _T_9260_11 : _T_12419; // @[Mux.scala 46:16:@10650.4]
  assign _T_12422 = 6'hb == _T_10211_35; // @[Mux.scala 46:19:@10651.4]
  assign _T_12423 = _T_12422 ? _T_9260_10 : _T_12421; // @[Mux.scala 46:16:@10652.4]
  assign _T_12424 = 6'ha == _T_10211_35; // @[Mux.scala 46:19:@10653.4]
  assign _T_12425 = _T_12424 ? _T_9260_9 : _T_12423; // @[Mux.scala 46:16:@10654.4]
  assign _T_12426 = 6'h9 == _T_10211_35; // @[Mux.scala 46:19:@10655.4]
  assign _T_12427 = _T_12426 ? _T_9260_8 : _T_12425; // @[Mux.scala 46:16:@10656.4]
  assign _T_12428 = 6'h8 == _T_10211_35; // @[Mux.scala 46:19:@10657.4]
  assign _T_12429 = _T_12428 ? _T_9260_7 : _T_12427; // @[Mux.scala 46:16:@10658.4]
  assign _T_12430 = 6'h7 == _T_10211_35; // @[Mux.scala 46:19:@10659.4]
  assign _T_12431 = _T_12430 ? _T_9260_6 : _T_12429; // @[Mux.scala 46:16:@10660.4]
  assign _T_12432 = 6'h6 == _T_10211_35; // @[Mux.scala 46:19:@10661.4]
  assign _T_12433 = _T_12432 ? _T_9260_5 : _T_12431; // @[Mux.scala 46:16:@10662.4]
  assign _T_12434 = 6'h5 == _T_10211_35; // @[Mux.scala 46:19:@10663.4]
  assign _T_12435 = _T_12434 ? _T_9260_4 : _T_12433; // @[Mux.scala 46:16:@10664.4]
  assign _T_12436 = 6'h4 == _T_10211_35; // @[Mux.scala 46:19:@10665.4]
  assign _T_12437 = _T_12436 ? _T_9260_3 : _T_12435; // @[Mux.scala 46:16:@10666.4]
  assign _T_12438 = 6'h3 == _T_10211_35; // @[Mux.scala 46:19:@10667.4]
  assign _T_12439 = _T_12438 ? _T_9260_2 : _T_12437; // @[Mux.scala 46:16:@10668.4]
  assign _T_12440 = 6'h2 == _T_10211_35; // @[Mux.scala 46:19:@10669.4]
  assign _T_12441 = _T_12440 ? _T_9260_1 : _T_12439; // @[Mux.scala 46:16:@10670.4]
  assign _T_12442 = 6'h1 == _T_10211_35; // @[Mux.scala 46:19:@10671.4]
  assign _T_12443 = _T_12442 ? _T_9260_0 : _T_12441; // @[Mux.scala 46:16:@10672.4]
  assign _T_12482 = 6'h25 == _T_10211_36; // @[Mux.scala 46:19:@10674.4]
  assign _T_12483 = _T_12482 ? _T_9260_36 : 8'h0; // @[Mux.scala 46:16:@10675.4]
  assign _T_12484 = 6'h24 == _T_10211_36; // @[Mux.scala 46:19:@10676.4]
  assign _T_12485 = _T_12484 ? _T_9260_35 : _T_12483; // @[Mux.scala 46:16:@10677.4]
  assign _T_12486 = 6'h23 == _T_10211_36; // @[Mux.scala 46:19:@10678.4]
  assign _T_12487 = _T_12486 ? _T_9260_34 : _T_12485; // @[Mux.scala 46:16:@10679.4]
  assign _T_12488 = 6'h22 == _T_10211_36; // @[Mux.scala 46:19:@10680.4]
  assign _T_12489 = _T_12488 ? _T_9260_33 : _T_12487; // @[Mux.scala 46:16:@10681.4]
  assign _T_12490 = 6'h21 == _T_10211_36; // @[Mux.scala 46:19:@10682.4]
  assign _T_12491 = _T_12490 ? _T_9260_32 : _T_12489; // @[Mux.scala 46:16:@10683.4]
  assign _T_12492 = 6'h20 == _T_10211_36; // @[Mux.scala 46:19:@10684.4]
  assign _T_12493 = _T_12492 ? _T_9260_31 : _T_12491; // @[Mux.scala 46:16:@10685.4]
  assign _T_12494 = 6'h1f == _T_10211_36; // @[Mux.scala 46:19:@10686.4]
  assign _T_12495 = _T_12494 ? _T_9260_30 : _T_12493; // @[Mux.scala 46:16:@10687.4]
  assign _T_12496 = 6'h1e == _T_10211_36; // @[Mux.scala 46:19:@10688.4]
  assign _T_12497 = _T_12496 ? _T_9260_29 : _T_12495; // @[Mux.scala 46:16:@10689.4]
  assign _T_12498 = 6'h1d == _T_10211_36; // @[Mux.scala 46:19:@10690.4]
  assign _T_12499 = _T_12498 ? _T_9260_28 : _T_12497; // @[Mux.scala 46:16:@10691.4]
  assign _T_12500 = 6'h1c == _T_10211_36; // @[Mux.scala 46:19:@10692.4]
  assign _T_12501 = _T_12500 ? _T_9260_27 : _T_12499; // @[Mux.scala 46:16:@10693.4]
  assign _T_12502 = 6'h1b == _T_10211_36; // @[Mux.scala 46:19:@10694.4]
  assign _T_12503 = _T_12502 ? _T_9260_26 : _T_12501; // @[Mux.scala 46:16:@10695.4]
  assign _T_12504 = 6'h1a == _T_10211_36; // @[Mux.scala 46:19:@10696.4]
  assign _T_12505 = _T_12504 ? _T_9260_25 : _T_12503; // @[Mux.scala 46:16:@10697.4]
  assign _T_12506 = 6'h19 == _T_10211_36; // @[Mux.scala 46:19:@10698.4]
  assign _T_12507 = _T_12506 ? _T_9260_24 : _T_12505; // @[Mux.scala 46:16:@10699.4]
  assign _T_12508 = 6'h18 == _T_10211_36; // @[Mux.scala 46:19:@10700.4]
  assign _T_12509 = _T_12508 ? _T_9260_23 : _T_12507; // @[Mux.scala 46:16:@10701.4]
  assign _T_12510 = 6'h17 == _T_10211_36; // @[Mux.scala 46:19:@10702.4]
  assign _T_12511 = _T_12510 ? _T_9260_22 : _T_12509; // @[Mux.scala 46:16:@10703.4]
  assign _T_12512 = 6'h16 == _T_10211_36; // @[Mux.scala 46:19:@10704.4]
  assign _T_12513 = _T_12512 ? _T_9260_21 : _T_12511; // @[Mux.scala 46:16:@10705.4]
  assign _T_12514 = 6'h15 == _T_10211_36; // @[Mux.scala 46:19:@10706.4]
  assign _T_12515 = _T_12514 ? _T_9260_20 : _T_12513; // @[Mux.scala 46:16:@10707.4]
  assign _T_12516 = 6'h14 == _T_10211_36; // @[Mux.scala 46:19:@10708.4]
  assign _T_12517 = _T_12516 ? _T_9260_19 : _T_12515; // @[Mux.scala 46:16:@10709.4]
  assign _T_12518 = 6'h13 == _T_10211_36; // @[Mux.scala 46:19:@10710.4]
  assign _T_12519 = _T_12518 ? _T_9260_18 : _T_12517; // @[Mux.scala 46:16:@10711.4]
  assign _T_12520 = 6'h12 == _T_10211_36; // @[Mux.scala 46:19:@10712.4]
  assign _T_12521 = _T_12520 ? _T_9260_17 : _T_12519; // @[Mux.scala 46:16:@10713.4]
  assign _T_12522 = 6'h11 == _T_10211_36; // @[Mux.scala 46:19:@10714.4]
  assign _T_12523 = _T_12522 ? _T_9260_16 : _T_12521; // @[Mux.scala 46:16:@10715.4]
  assign _T_12524 = 6'h10 == _T_10211_36; // @[Mux.scala 46:19:@10716.4]
  assign _T_12525 = _T_12524 ? _T_9260_15 : _T_12523; // @[Mux.scala 46:16:@10717.4]
  assign _T_12526 = 6'hf == _T_10211_36; // @[Mux.scala 46:19:@10718.4]
  assign _T_12527 = _T_12526 ? _T_9260_14 : _T_12525; // @[Mux.scala 46:16:@10719.4]
  assign _T_12528 = 6'he == _T_10211_36; // @[Mux.scala 46:19:@10720.4]
  assign _T_12529 = _T_12528 ? _T_9260_13 : _T_12527; // @[Mux.scala 46:16:@10721.4]
  assign _T_12530 = 6'hd == _T_10211_36; // @[Mux.scala 46:19:@10722.4]
  assign _T_12531 = _T_12530 ? _T_9260_12 : _T_12529; // @[Mux.scala 46:16:@10723.4]
  assign _T_12532 = 6'hc == _T_10211_36; // @[Mux.scala 46:19:@10724.4]
  assign _T_12533 = _T_12532 ? _T_9260_11 : _T_12531; // @[Mux.scala 46:16:@10725.4]
  assign _T_12534 = 6'hb == _T_10211_36; // @[Mux.scala 46:19:@10726.4]
  assign _T_12535 = _T_12534 ? _T_9260_10 : _T_12533; // @[Mux.scala 46:16:@10727.4]
  assign _T_12536 = 6'ha == _T_10211_36; // @[Mux.scala 46:19:@10728.4]
  assign _T_12537 = _T_12536 ? _T_9260_9 : _T_12535; // @[Mux.scala 46:16:@10729.4]
  assign _T_12538 = 6'h9 == _T_10211_36; // @[Mux.scala 46:19:@10730.4]
  assign _T_12539 = _T_12538 ? _T_9260_8 : _T_12537; // @[Mux.scala 46:16:@10731.4]
  assign _T_12540 = 6'h8 == _T_10211_36; // @[Mux.scala 46:19:@10732.4]
  assign _T_12541 = _T_12540 ? _T_9260_7 : _T_12539; // @[Mux.scala 46:16:@10733.4]
  assign _T_12542 = 6'h7 == _T_10211_36; // @[Mux.scala 46:19:@10734.4]
  assign _T_12543 = _T_12542 ? _T_9260_6 : _T_12541; // @[Mux.scala 46:16:@10735.4]
  assign _T_12544 = 6'h6 == _T_10211_36; // @[Mux.scala 46:19:@10736.4]
  assign _T_12545 = _T_12544 ? _T_9260_5 : _T_12543; // @[Mux.scala 46:16:@10737.4]
  assign _T_12546 = 6'h5 == _T_10211_36; // @[Mux.scala 46:19:@10738.4]
  assign _T_12547 = _T_12546 ? _T_9260_4 : _T_12545; // @[Mux.scala 46:16:@10739.4]
  assign _T_12548 = 6'h4 == _T_10211_36; // @[Mux.scala 46:19:@10740.4]
  assign _T_12549 = _T_12548 ? _T_9260_3 : _T_12547; // @[Mux.scala 46:16:@10741.4]
  assign _T_12550 = 6'h3 == _T_10211_36; // @[Mux.scala 46:19:@10742.4]
  assign _T_12551 = _T_12550 ? _T_9260_2 : _T_12549; // @[Mux.scala 46:16:@10743.4]
  assign _T_12552 = 6'h2 == _T_10211_36; // @[Mux.scala 46:19:@10744.4]
  assign _T_12553 = _T_12552 ? _T_9260_1 : _T_12551; // @[Mux.scala 46:16:@10745.4]
  assign _T_12554 = 6'h1 == _T_10211_36; // @[Mux.scala 46:19:@10746.4]
  assign _T_12555 = _T_12554 ? _T_9260_0 : _T_12553; // @[Mux.scala 46:16:@10747.4]
  assign _T_12595 = 6'h26 == _T_10211_37; // @[Mux.scala 46:19:@10749.4]
  assign _T_12596 = _T_12595 ? _T_9260_37 : 8'h0; // @[Mux.scala 46:16:@10750.4]
  assign _T_12597 = 6'h25 == _T_10211_37; // @[Mux.scala 46:19:@10751.4]
  assign _T_12598 = _T_12597 ? _T_9260_36 : _T_12596; // @[Mux.scala 46:16:@10752.4]
  assign _T_12599 = 6'h24 == _T_10211_37; // @[Mux.scala 46:19:@10753.4]
  assign _T_12600 = _T_12599 ? _T_9260_35 : _T_12598; // @[Mux.scala 46:16:@10754.4]
  assign _T_12601 = 6'h23 == _T_10211_37; // @[Mux.scala 46:19:@10755.4]
  assign _T_12602 = _T_12601 ? _T_9260_34 : _T_12600; // @[Mux.scala 46:16:@10756.4]
  assign _T_12603 = 6'h22 == _T_10211_37; // @[Mux.scala 46:19:@10757.4]
  assign _T_12604 = _T_12603 ? _T_9260_33 : _T_12602; // @[Mux.scala 46:16:@10758.4]
  assign _T_12605 = 6'h21 == _T_10211_37; // @[Mux.scala 46:19:@10759.4]
  assign _T_12606 = _T_12605 ? _T_9260_32 : _T_12604; // @[Mux.scala 46:16:@10760.4]
  assign _T_12607 = 6'h20 == _T_10211_37; // @[Mux.scala 46:19:@10761.4]
  assign _T_12608 = _T_12607 ? _T_9260_31 : _T_12606; // @[Mux.scala 46:16:@10762.4]
  assign _T_12609 = 6'h1f == _T_10211_37; // @[Mux.scala 46:19:@10763.4]
  assign _T_12610 = _T_12609 ? _T_9260_30 : _T_12608; // @[Mux.scala 46:16:@10764.4]
  assign _T_12611 = 6'h1e == _T_10211_37; // @[Mux.scala 46:19:@10765.4]
  assign _T_12612 = _T_12611 ? _T_9260_29 : _T_12610; // @[Mux.scala 46:16:@10766.4]
  assign _T_12613 = 6'h1d == _T_10211_37; // @[Mux.scala 46:19:@10767.4]
  assign _T_12614 = _T_12613 ? _T_9260_28 : _T_12612; // @[Mux.scala 46:16:@10768.4]
  assign _T_12615 = 6'h1c == _T_10211_37; // @[Mux.scala 46:19:@10769.4]
  assign _T_12616 = _T_12615 ? _T_9260_27 : _T_12614; // @[Mux.scala 46:16:@10770.4]
  assign _T_12617 = 6'h1b == _T_10211_37; // @[Mux.scala 46:19:@10771.4]
  assign _T_12618 = _T_12617 ? _T_9260_26 : _T_12616; // @[Mux.scala 46:16:@10772.4]
  assign _T_12619 = 6'h1a == _T_10211_37; // @[Mux.scala 46:19:@10773.4]
  assign _T_12620 = _T_12619 ? _T_9260_25 : _T_12618; // @[Mux.scala 46:16:@10774.4]
  assign _T_12621 = 6'h19 == _T_10211_37; // @[Mux.scala 46:19:@10775.4]
  assign _T_12622 = _T_12621 ? _T_9260_24 : _T_12620; // @[Mux.scala 46:16:@10776.4]
  assign _T_12623 = 6'h18 == _T_10211_37; // @[Mux.scala 46:19:@10777.4]
  assign _T_12624 = _T_12623 ? _T_9260_23 : _T_12622; // @[Mux.scala 46:16:@10778.4]
  assign _T_12625 = 6'h17 == _T_10211_37; // @[Mux.scala 46:19:@10779.4]
  assign _T_12626 = _T_12625 ? _T_9260_22 : _T_12624; // @[Mux.scala 46:16:@10780.4]
  assign _T_12627 = 6'h16 == _T_10211_37; // @[Mux.scala 46:19:@10781.4]
  assign _T_12628 = _T_12627 ? _T_9260_21 : _T_12626; // @[Mux.scala 46:16:@10782.4]
  assign _T_12629 = 6'h15 == _T_10211_37; // @[Mux.scala 46:19:@10783.4]
  assign _T_12630 = _T_12629 ? _T_9260_20 : _T_12628; // @[Mux.scala 46:16:@10784.4]
  assign _T_12631 = 6'h14 == _T_10211_37; // @[Mux.scala 46:19:@10785.4]
  assign _T_12632 = _T_12631 ? _T_9260_19 : _T_12630; // @[Mux.scala 46:16:@10786.4]
  assign _T_12633 = 6'h13 == _T_10211_37; // @[Mux.scala 46:19:@10787.4]
  assign _T_12634 = _T_12633 ? _T_9260_18 : _T_12632; // @[Mux.scala 46:16:@10788.4]
  assign _T_12635 = 6'h12 == _T_10211_37; // @[Mux.scala 46:19:@10789.4]
  assign _T_12636 = _T_12635 ? _T_9260_17 : _T_12634; // @[Mux.scala 46:16:@10790.4]
  assign _T_12637 = 6'h11 == _T_10211_37; // @[Mux.scala 46:19:@10791.4]
  assign _T_12638 = _T_12637 ? _T_9260_16 : _T_12636; // @[Mux.scala 46:16:@10792.4]
  assign _T_12639 = 6'h10 == _T_10211_37; // @[Mux.scala 46:19:@10793.4]
  assign _T_12640 = _T_12639 ? _T_9260_15 : _T_12638; // @[Mux.scala 46:16:@10794.4]
  assign _T_12641 = 6'hf == _T_10211_37; // @[Mux.scala 46:19:@10795.4]
  assign _T_12642 = _T_12641 ? _T_9260_14 : _T_12640; // @[Mux.scala 46:16:@10796.4]
  assign _T_12643 = 6'he == _T_10211_37; // @[Mux.scala 46:19:@10797.4]
  assign _T_12644 = _T_12643 ? _T_9260_13 : _T_12642; // @[Mux.scala 46:16:@10798.4]
  assign _T_12645 = 6'hd == _T_10211_37; // @[Mux.scala 46:19:@10799.4]
  assign _T_12646 = _T_12645 ? _T_9260_12 : _T_12644; // @[Mux.scala 46:16:@10800.4]
  assign _T_12647 = 6'hc == _T_10211_37; // @[Mux.scala 46:19:@10801.4]
  assign _T_12648 = _T_12647 ? _T_9260_11 : _T_12646; // @[Mux.scala 46:16:@10802.4]
  assign _T_12649 = 6'hb == _T_10211_37; // @[Mux.scala 46:19:@10803.4]
  assign _T_12650 = _T_12649 ? _T_9260_10 : _T_12648; // @[Mux.scala 46:16:@10804.4]
  assign _T_12651 = 6'ha == _T_10211_37; // @[Mux.scala 46:19:@10805.4]
  assign _T_12652 = _T_12651 ? _T_9260_9 : _T_12650; // @[Mux.scala 46:16:@10806.4]
  assign _T_12653 = 6'h9 == _T_10211_37; // @[Mux.scala 46:19:@10807.4]
  assign _T_12654 = _T_12653 ? _T_9260_8 : _T_12652; // @[Mux.scala 46:16:@10808.4]
  assign _T_12655 = 6'h8 == _T_10211_37; // @[Mux.scala 46:19:@10809.4]
  assign _T_12656 = _T_12655 ? _T_9260_7 : _T_12654; // @[Mux.scala 46:16:@10810.4]
  assign _T_12657 = 6'h7 == _T_10211_37; // @[Mux.scala 46:19:@10811.4]
  assign _T_12658 = _T_12657 ? _T_9260_6 : _T_12656; // @[Mux.scala 46:16:@10812.4]
  assign _T_12659 = 6'h6 == _T_10211_37; // @[Mux.scala 46:19:@10813.4]
  assign _T_12660 = _T_12659 ? _T_9260_5 : _T_12658; // @[Mux.scala 46:16:@10814.4]
  assign _T_12661 = 6'h5 == _T_10211_37; // @[Mux.scala 46:19:@10815.4]
  assign _T_12662 = _T_12661 ? _T_9260_4 : _T_12660; // @[Mux.scala 46:16:@10816.4]
  assign _T_12663 = 6'h4 == _T_10211_37; // @[Mux.scala 46:19:@10817.4]
  assign _T_12664 = _T_12663 ? _T_9260_3 : _T_12662; // @[Mux.scala 46:16:@10818.4]
  assign _T_12665 = 6'h3 == _T_10211_37; // @[Mux.scala 46:19:@10819.4]
  assign _T_12666 = _T_12665 ? _T_9260_2 : _T_12664; // @[Mux.scala 46:16:@10820.4]
  assign _T_12667 = 6'h2 == _T_10211_37; // @[Mux.scala 46:19:@10821.4]
  assign _T_12668 = _T_12667 ? _T_9260_1 : _T_12666; // @[Mux.scala 46:16:@10822.4]
  assign _T_12669 = 6'h1 == _T_10211_37; // @[Mux.scala 46:19:@10823.4]
  assign _T_12670 = _T_12669 ? _T_9260_0 : _T_12668; // @[Mux.scala 46:16:@10824.4]
  assign _T_12711 = 6'h27 == _T_10211_38; // @[Mux.scala 46:19:@10826.4]
  assign _T_12712 = _T_12711 ? _T_9260_38 : 8'h0; // @[Mux.scala 46:16:@10827.4]
  assign _T_12713 = 6'h26 == _T_10211_38; // @[Mux.scala 46:19:@10828.4]
  assign _T_12714 = _T_12713 ? _T_9260_37 : _T_12712; // @[Mux.scala 46:16:@10829.4]
  assign _T_12715 = 6'h25 == _T_10211_38; // @[Mux.scala 46:19:@10830.4]
  assign _T_12716 = _T_12715 ? _T_9260_36 : _T_12714; // @[Mux.scala 46:16:@10831.4]
  assign _T_12717 = 6'h24 == _T_10211_38; // @[Mux.scala 46:19:@10832.4]
  assign _T_12718 = _T_12717 ? _T_9260_35 : _T_12716; // @[Mux.scala 46:16:@10833.4]
  assign _T_12719 = 6'h23 == _T_10211_38; // @[Mux.scala 46:19:@10834.4]
  assign _T_12720 = _T_12719 ? _T_9260_34 : _T_12718; // @[Mux.scala 46:16:@10835.4]
  assign _T_12721 = 6'h22 == _T_10211_38; // @[Mux.scala 46:19:@10836.4]
  assign _T_12722 = _T_12721 ? _T_9260_33 : _T_12720; // @[Mux.scala 46:16:@10837.4]
  assign _T_12723 = 6'h21 == _T_10211_38; // @[Mux.scala 46:19:@10838.4]
  assign _T_12724 = _T_12723 ? _T_9260_32 : _T_12722; // @[Mux.scala 46:16:@10839.4]
  assign _T_12725 = 6'h20 == _T_10211_38; // @[Mux.scala 46:19:@10840.4]
  assign _T_12726 = _T_12725 ? _T_9260_31 : _T_12724; // @[Mux.scala 46:16:@10841.4]
  assign _T_12727 = 6'h1f == _T_10211_38; // @[Mux.scala 46:19:@10842.4]
  assign _T_12728 = _T_12727 ? _T_9260_30 : _T_12726; // @[Mux.scala 46:16:@10843.4]
  assign _T_12729 = 6'h1e == _T_10211_38; // @[Mux.scala 46:19:@10844.4]
  assign _T_12730 = _T_12729 ? _T_9260_29 : _T_12728; // @[Mux.scala 46:16:@10845.4]
  assign _T_12731 = 6'h1d == _T_10211_38; // @[Mux.scala 46:19:@10846.4]
  assign _T_12732 = _T_12731 ? _T_9260_28 : _T_12730; // @[Mux.scala 46:16:@10847.4]
  assign _T_12733 = 6'h1c == _T_10211_38; // @[Mux.scala 46:19:@10848.4]
  assign _T_12734 = _T_12733 ? _T_9260_27 : _T_12732; // @[Mux.scala 46:16:@10849.4]
  assign _T_12735 = 6'h1b == _T_10211_38; // @[Mux.scala 46:19:@10850.4]
  assign _T_12736 = _T_12735 ? _T_9260_26 : _T_12734; // @[Mux.scala 46:16:@10851.4]
  assign _T_12737 = 6'h1a == _T_10211_38; // @[Mux.scala 46:19:@10852.4]
  assign _T_12738 = _T_12737 ? _T_9260_25 : _T_12736; // @[Mux.scala 46:16:@10853.4]
  assign _T_12739 = 6'h19 == _T_10211_38; // @[Mux.scala 46:19:@10854.4]
  assign _T_12740 = _T_12739 ? _T_9260_24 : _T_12738; // @[Mux.scala 46:16:@10855.4]
  assign _T_12741 = 6'h18 == _T_10211_38; // @[Mux.scala 46:19:@10856.4]
  assign _T_12742 = _T_12741 ? _T_9260_23 : _T_12740; // @[Mux.scala 46:16:@10857.4]
  assign _T_12743 = 6'h17 == _T_10211_38; // @[Mux.scala 46:19:@10858.4]
  assign _T_12744 = _T_12743 ? _T_9260_22 : _T_12742; // @[Mux.scala 46:16:@10859.4]
  assign _T_12745 = 6'h16 == _T_10211_38; // @[Mux.scala 46:19:@10860.4]
  assign _T_12746 = _T_12745 ? _T_9260_21 : _T_12744; // @[Mux.scala 46:16:@10861.4]
  assign _T_12747 = 6'h15 == _T_10211_38; // @[Mux.scala 46:19:@10862.4]
  assign _T_12748 = _T_12747 ? _T_9260_20 : _T_12746; // @[Mux.scala 46:16:@10863.4]
  assign _T_12749 = 6'h14 == _T_10211_38; // @[Mux.scala 46:19:@10864.4]
  assign _T_12750 = _T_12749 ? _T_9260_19 : _T_12748; // @[Mux.scala 46:16:@10865.4]
  assign _T_12751 = 6'h13 == _T_10211_38; // @[Mux.scala 46:19:@10866.4]
  assign _T_12752 = _T_12751 ? _T_9260_18 : _T_12750; // @[Mux.scala 46:16:@10867.4]
  assign _T_12753 = 6'h12 == _T_10211_38; // @[Mux.scala 46:19:@10868.4]
  assign _T_12754 = _T_12753 ? _T_9260_17 : _T_12752; // @[Mux.scala 46:16:@10869.4]
  assign _T_12755 = 6'h11 == _T_10211_38; // @[Mux.scala 46:19:@10870.4]
  assign _T_12756 = _T_12755 ? _T_9260_16 : _T_12754; // @[Mux.scala 46:16:@10871.4]
  assign _T_12757 = 6'h10 == _T_10211_38; // @[Mux.scala 46:19:@10872.4]
  assign _T_12758 = _T_12757 ? _T_9260_15 : _T_12756; // @[Mux.scala 46:16:@10873.4]
  assign _T_12759 = 6'hf == _T_10211_38; // @[Mux.scala 46:19:@10874.4]
  assign _T_12760 = _T_12759 ? _T_9260_14 : _T_12758; // @[Mux.scala 46:16:@10875.4]
  assign _T_12761 = 6'he == _T_10211_38; // @[Mux.scala 46:19:@10876.4]
  assign _T_12762 = _T_12761 ? _T_9260_13 : _T_12760; // @[Mux.scala 46:16:@10877.4]
  assign _T_12763 = 6'hd == _T_10211_38; // @[Mux.scala 46:19:@10878.4]
  assign _T_12764 = _T_12763 ? _T_9260_12 : _T_12762; // @[Mux.scala 46:16:@10879.4]
  assign _T_12765 = 6'hc == _T_10211_38; // @[Mux.scala 46:19:@10880.4]
  assign _T_12766 = _T_12765 ? _T_9260_11 : _T_12764; // @[Mux.scala 46:16:@10881.4]
  assign _T_12767 = 6'hb == _T_10211_38; // @[Mux.scala 46:19:@10882.4]
  assign _T_12768 = _T_12767 ? _T_9260_10 : _T_12766; // @[Mux.scala 46:16:@10883.4]
  assign _T_12769 = 6'ha == _T_10211_38; // @[Mux.scala 46:19:@10884.4]
  assign _T_12770 = _T_12769 ? _T_9260_9 : _T_12768; // @[Mux.scala 46:16:@10885.4]
  assign _T_12771 = 6'h9 == _T_10211_38; // @[Mux.scala 46:19:@10886.4]
  assign _T_12772 = _T_12771 ? _T_9260_8 : _T_12770; // @[Mux.scala 46:16:@10887.4]
  assign _T_12773 = 6'h8 == _T_10211_38; // @[Mux.scala 46:19:@10888.4]
  assign _T_12774 = _T_12773 ? _T_9260_7 : _T_12772; // @[Mux.scala 46:16:@10889.4]
  assign _T_12775 = 6'h7 == _T_10211_38; // @[Mux.scala 46:19:@10890.4]
  assign _T_12776 = _T_12775 ? _T_9260_6 : _T_12774; // @[Mux.scala 46:16:@10891.4]
  assign _T_12777 = 6'h6 == _T_10211_38; // @[Mux.scala 46:19:@10892.4]
  assign _T_12778 = _T_12777 ? _T_9260_5 : _T_12776; // @[Mux.scala 46:16:@10893.4]
  assign _T_12779 = 6'h5 == _T_10211_38; // @[Mux.scala 46:19:@10894.4]
  assign _T_12780 = _T_12779 ? _T_9260_4 : _T_12778; // @[Mux.scala 46:16:@10895.4]
  assign _T_12781 = 6'h4 == _T_10211_38; // @[Mux.scala 46:19:@10896.4]
  assign _T_12782 = _T_12781 ? _T_9260_3 : _T_12780; // @[Mux.scala 46:16:@10897.4]
  assign _T_12783 = 6'h3 == _T_10211_38; // @[Mux.scala 46:19:@10898.4]
  assign _T_12784 = _T_12783 ? _T_9260_2 : _T_12782; // @[Mux.scala 46:16:@10899.4]
  assign _T_12785 = 6'h2 == _T_10211_38; // @[Mux.scala 46:19:@10900.4]
  assign _T_12786 = _T_12785 ? _T_9260_1 : _T_12784; // @[Mux.scala 46:16:@10901.4]
  assign _T_12787 = 6'h1 == _T_10211_38; // @[Mux.scala 46:19:@10902.4]
  assign _T_12788 = _T_12787 ? _T_9260_0 : _T_12786; // @[Mux.scala 46:16:@10903.4]
  assign _T_12830 = 6'h28 == _T_10211_39; // @[Mux.scala 46:19:@10905.4]
  assign _T_12831 = _T_12830 ? _T_9260_39 : 8'h0; // @[Mux.scala 46:16:@10906.4]
  assign _T_12832 = 6'h27 == _T_10211_39; // @[Mux.scala 46:19:@10907.4]
  assign _T_12833 = _T_12832 ? _T_9260_38 : _T_12831; // @[Mux.scala 46:16:@10908.4]
  assign _T_12834 = 6'h26 == _T_10211_39; // @[Mux.scala 46:19:@10909.4]
  assign _T_12835 = _T_12834 ? _T_9260_37 : _T_12833; // @[Mux.scala 46:16:@10910.4]
  assign _T_12836 = 6'h25 == _T_10211_39; // @[Mux.scala 46:19:@10911.4]
  assign _T_12837 = _T_12836 ? _T_9260_36 : _T_12835; // @[Mux.scala 46:16:@10912.4]
  assign _T_12838 = 6'h24 == _T_10211_39; // @[Mux.scala 46:19:@10913.4]
  assign _T_12839 = _T_12838 ? _T_9260_35 : _T_12837; // @[Mux.scala 46:16:@10914.4]
  assign _T_12840 = 6'h23 == _T_10211_39; // @[Mux.scala 46:19:@10915.4]
  assign _T_12841 = _T_12840 ? _T_9260_34 : _T_12839; // @[Mux.scala 46:16:@10916.4]
  assign _T_12842 = 6'h22 == _T_10211_39; // @[Mux.scala 46:19:@10917.4]
  assign _T_12843 = _T_12842 ? _T_9260_33 : _T_12841; // @[Mux.scala 46:16:@10918.4]
  assign _T_12844 = 6'h21 == _T_10211_39; // @[Mux.scala 46:19:@10919.4]
  assign _T_12845 = _T_12844 ? _T_9260_32 : _T_12843; // @[Mux.scala 46:16:@10920.4]
  assign _T_12846 = 6'h20 == _T_10211_39; // @[Mux.scala 46:19:@10921.4]
  assign _T_12847 = _T_12846 ? _T_9260_31 : _T_12845; // @[Mux.scala 46:16:@10922.4]
  assign _T_12848 = 6'h1f == _T_10211_39; // @[Mux.scala 46:19:@10923.4]
  assign _T_12849 = _T_12848 ? _T_9260_30 : _T_12847; // @[Mux.scala 46:16:@10924.4]
  assign _T_12850 = 6'h1e == _T_10211_39; // @[Mux.scala 46:19:@10925.4]
  assign _T_12851 = _T_12850 ? _T_9260_29 : _T_12849; // @[Mux.scala 46:16:@10926.4]
  assign _T_12852 = 6'h1d == _T_10211_39; // @[Mux.scala 46:19:@10927.4]
  assign _T_12853 = _T_12852 ? _T_9260_28 : _T_12851; // @[Mux.scala 46:16:@10928.4]
  assign _T_12854 = 6'h1c == _T_10211_39; // @[Mux.scala 46:19:@10929.4]
  assign _T_12855 = _T_12854 ? _T_9260_27 : _T_12853; // @[Mux.scala 46:16:@10930.4]
  assign _T_12856 = 6'h1b == _T_10211_39; // @[Mux.scala 46:19:@10931.4]
  assign _T_12857 = _T_12856 ? _T_9260_26 : _T_12855; // @[Mux.scala 46:16:@10932.4]
  assign _T_12858 = 6'h1a == _T_10211_39; // @[Mux.scala 46:19:@10933.4]
  assign _T_12859 = _T_12858 ? _T_9260_25 : _T_12857; // @[Mux.scala 46:16:@10934.4]
  assign _T_12860 = 6'h19 == _T_10211_39; // @[Mux.scala 46:19:@10935.4]
  assign _T_12861 = _T_12860 ? _T_9260_24 : _T_12859; // @[Mux.scala 46:16:@10936.4]
  assign _T_12862 = 6'h18 == _T_10211_39; // @[Mux.scala 46:19:@10937.4]
  assign _T_12863 = _T_12862 ? _T_9260_23 : _T_12861; // @[Mux.scala 46:16:@10938.4]
  assign _T_12864 = 6'h17 == _T_10211_39; // @[Mux.scala 46:19:@10939.4]
  assign _T_12865 = _T_12864 ? _T_9260_22 : _T_12863; // @[Mux.scala 46:16:@10940.4]
  assign _T_12866 = 6'h16 == _T_10211_39; // @[Mux.scala 46:19:@10941.4]
  assign _T_12867 = _T_12866 ? _T_9260_21 : _T_12865; // @[Mux.scala 46:16:@10942.4]
  assign _T_12868 = 6'h15 == _T_10211_39; // @[Mux.scala 46:19:@10943.4]
  assign _T_12869 = _T_12868 ? _T_9260_20 : _T_12867; // @[Mux.scala 46:16:@10944.4]
  assign _T_12870 = 6'h14 == _T_10211_39; // @[Mux.scala 46:19:@10945.4]
  assign _T_12871 = _T_12870 ? _T_9260_19 : _T_12869; // @[Mux.scala 46:16:@10946.4]
  assign _T_12872 = 6'h13 == _T_10211_39; // @[Mux.scala 46:19:@10947.4]
  assign _T_12873 = _T_12872 ? _T_9260_18 : _T_12871; // @[Mux.scala 46:16:@10948.4]
  assign _T_12874 = 6'h12 == _T_10211_39; // @[Mux.scala 46:19:@10949.4]
  assign _T_12875 = _T_12874 ? _T_9260_17 : _T_12873; // @[Mux.scala 46:16:@10950.4]
  assign _T_12876 = 6'h11 == _T_10211_39; // @[Mux.scala 46:19:@10951.4]
  assign _T_12877 = _T_12876 ? _T_9260_16 : _T_12875; // @[Mux.scala 46:16:@10952.4]
  assign _T_12878 = 6'h10 == _T_10211_39; // @[Mux.scala 46:19:@10953.4]
  assign _T_12879 = _T_12878 ? _T_9260_15 : _T_12877; // @[Mux.scala 46:16:@10954.4]
  assign _T_12880 = 6'hf == _T_10211_39; // @[Mux.scala 46:19:@10955.4]
  assign _T_12881 = _T_12880 ? _T_9260_14 : _T_12879; // @[Mux.scala 46:16:@10956.4]
  assign _T_12882 = 6'he == _T_10211_39; // @[Mux.scala 46:19:@10957.4]
  assign _T_12883 = _T_12882 ? _T_9260_13 : _T_12881; // @[Mux.scala 46:16:@10958.4]
  assign _T_12884 = 6'hd == _T_10211_39; // @[Mux.scala 46:19:@10959.4]
  assign _T_12885 = _T_12884 ? _T_9260_12 : _T_12883; // @[Mux.scala 46:16:@10960.4]
  assign _T_12886 = 6'hc == _T_10211_39; // @[Mux.scala 46:19:@10961.4]
  assign _T_12887 = _T_12886 ? _T_9260_11 : _T_12885; // @[Mux.scala 46:16:@10962.4]
  assign _T_12888 = 6'hb == _T_10211_39; // @[Mux.scala 46:19:@10963.4]
  assign _T_12889 = _T_12888 ? _T_9260_10 : _T_12887; // @[Mux.scala 46:16:@10964.4]
  assign _T_12890 = 6'ha == _T_10211_39; // @[Mux.scala 46:19:@10965.4]
  assign _T_12891 = _T_12890 ? _T_9260_9 : _T_12889; // @[Mux.scala 46:16:@10966.4]
  assign _T_12892 = 6'h9 == _T_10211_39; // @[Mux.scala 46:19:@10967.4]
  assign _T_12893 = _T_12892 ? _T_9260_8 : _T_12891; // @[Mux.scala 46:16:@10968.4]
  assign _T_12894 = 6'h8 == _T_10211_39; // @[Mux.scala 46:19:@10969.4]
  assign _T_12895 = _T_12894 ? _T_9260_7 : _T_12893; // @[Mux.scala 46:16:@10970.4]
  assign _T_12896 = 6'h7 == _T_10211_39; // @[Mux.scala 46:19:@10971.4]
  assign _T_12897 = _T_12896 ? _T_9260_6 : _T_12895; // @[Mux.scala 46:16:@10972.4]
  assign _T_12898 = 6'h6 == _T_10211_39; // @[Mux.scala 46:19:@10973.4]
  assign _T_12899 = _T_12898 ? _T_9260_5 : _T_12897; // @[Mux.scala 46:16:@10974.4]
  assign _T_12900 = 6'h5 == _T_10211_39; // @[Mux.scala 46:19:@10975.4]
  assign _T_12901 = _T_12900 ? _T_9260_4 : _T_12899; // @[Mux.scala 46:16:@10976.4]
  assign _T_12902 = 6'h4 == _T_10211_39; // @[Mux.scala 46:19:@10977.4]
  assign _T_12903 = _T_12902 ? _T_9260_3 : _T_12901; // @[Mux.scala 46:16:@10978.4]
  assign _T_12904 = 6'h3 == _T_10211_39; // @[Mux.scala 46:19:@10979.4]
  assign _T_12905 = _T_12904 ? _T_9260_2 : _T_12903; // @[Mux.scala 46:16:@10980.4]
  assign _T_12906 = 6'h2 == _T_10211_39; // @[Mux.scala 46:19:@10981.4]
  assign _T_12907 = _T_12906 ? _T_9260_1 : _T_12905; // @[Mux.scala 46:16:@10982.4]
  assign _T_12908 = 6'h1 == _T_10211_39; // @[Mux.scala 46:19:@10983.4]
  assign _T_12909 = _T_12908 ? _T_9260_0 : _T_12907; // @[Mux.scala 46:16:@10984.4]
  assign _T_12952 = 6'h29 == _T_10211_40; // @[Mux.scala 46:19:@10986.4]
  assign _T_12953 = _T_12952 ? _T_9260_40 : 8'h0; // @[Mux.scala 46:16:@10987.4]
  assign _T_12954 = 6'h28 == _T_10211_40; // @[Mux.scala 46:19:@10988.4]
  assign _T_12955 = _T_12954 ? _T_9260_39 : _T_12953; // @[Mux.scala 46:16:@10989.4]
  assign _T_12956 = 6'h27 == _T_10211_40; // @[Mux.scala 46:19:@10990.4]
  assign _T_12957 = _T_12956 ? _T_9260_38 : _T_12955; // @[Mux.scala 46:16:@10991.4]
  assign _T_12958 = 6'h26 == _T_10211_40; // @[Mux.scala 46:19:@10992.4]
  assign _T_12959 = _T_12958 ? _T_9260_37 : _T_12957; // @[Mux.scala 46:16:@10993.4]
  assign _T_12960 = 6'h25 == _T_10211_40; // @[Mux.scala 46:19:@10994.4]
  assign _T_12961 = _T_12960 ? _T_9260_36 : _T_12959; // @[Mux.scala 46:16:@10995.4]
  assign _T_12962 = 6'h24 == _T_10211_40; // @[Mux.scala 46:19:@10996.4]
  assign _T_12963 = _T_12962 ? _T_9260_35 : _T_12961; // @[Mux.scala 46:16:@10997.4]
  assign _T_12964 = 6'h23 == _T_10211_40; // @[Mux.scala 46:19:@10998.4]
  assign _T_12965 = _T_12964 ? _T_9260_34 : _T_12963; // @[Mux.scala 46:16:@10999.4]
  assign _T_12966 = 6'h22 == _T_10211_40; // @[Mux.scala 46:19:@11000.4]
  assign _T_12967 = _T_12966 ? _T_9260_33 : _T_12965; // @[Mux.scala 46:16:@11001.4]
  assign _T_12968 = 6'h21 == _T_10211_40; // @[Mux.scala 46:19:@11002.4]
  assign _T_12969 = _T_12968 ? _T_9260_32 : _T_12967; // @[Mux.scala 46:16:@11003.4]
  assign _T_12970 = 6'h20 == _T_10211_40; // @[Mux.scala 46:19:@11004.4]
  assign _T_12971 = _T_12970 ? _T_9260_31 : _T_12969; // @[Mux.scala 46:16:@11005.4]
  assign _T_12972 = 6'h1f == _T_10211_40; // @[Mux.scala 46:19:@11006.4]
  assign _T_12973 = _T_12972 ? _T_9260_30 : _T_12971; // @[Mux.scala 46:16:@11007.4]
  assign _T_12974 = 6'h1e == _T_10211_40; // @[Mux.scala 46:19:@11008.4]
  assign _T_12975 = _T_12974 ? _T_9260_29 : _T_12973; // @[Mux.scala 46:16:@11009.4]
  assign _T_12976 = 6'h1d == _T_10211_40; // @[Mux.scala 46:19:@11010.4]
  assign _T_12977 = _T_12976 ? _T_9260_28 : _T_12975; // @[Mux.scala 46:16:@11011.4]
  assign _T_12978 = 6'h1c == _T_10211_40; // @[Mux.scala 46:19:@11012.4]
  assign _T_12979 = _T_12978 ? _T_9260_27 : _T_12977; // @[Mux.scala 46:16:@11013.4]
  assign _T_12980 = 6'h1b == _T_10211_40; // @[Mux.scala 46:19:@11014.4]
  assign _T_12981 = _T_12980 ? _T_9260_26 : _T_12979; // @[Mux.scala 46:16:@11015.4]
  assign _T_12982 = 6'h1a == _T_10211_40; // @[Mux.scala 46:19:@11016.4]
  assign _T_12983 = _T_12982 ? _T_9260_25 : _T_12981; // @[Mux.scala 46:16:@11017.4]
  assign _T_12984 = 6'h19 == _T_10211_40; // @[Mux.scala 46:19:@11018.4]
  assign _T_12985 = _T_12984 ? _T_9260_24 : _T_12983; // @[Mux.scala 46:16:@11019.4]
  assign _T_12986 = 6'h18 == _T_10211_40; // @[Mux.scala 46:19:@11020.4]
  assign _T_12987 = _T_12986 ? _T_9260_23 : _T_12985; // @[Mux.scala 46:16:@11021.4]
  assign _T_12988 = 6'h17 == _T_10211_40; // @[Mux.scala 46:19:@11022.4]
  assign _T_12989 = _T_12988 ? _T_9260_22 : _T_12987; // @[Mux.scala 46:16:@11023.4]
  assign _T_12990 = 6'h16 == _T_10211_40; // @[Mux.scala 46:19:@11024.4]
  assign _T_12991 = _T_12990 ? _T_9260_21 : _T_12989; // @[Mux.scala 46:16:@11025.4]
  assign _T_12992 = 6'h15 == _T_10211_40; // @[Mux.scala 46:19:@11026.4]
  assign _T_12993 = _T_12992 ? _T_9260_20 : _T_12991; // @[Mux.scala 46:16:@11027.4]
  assign _T_12994 = 6'h14 == _T_10211_40; // @[Mux.scala 46:19:@11028.4]
  assign _T_12995 = _T_12994 ? _T_9260_19 : _T_12993; // @[Mux.scala 46:16:@11029.4]
  assign _T_12996 = 6'h13 == _T_10211_40; // @[Mux.scala 46:19:@11030.4]
  assign _T_12997 = _T_12996 ? _T_9260_18 : _T_12995; // @[Mux.scala 46:16:@11031.4]
  assign _T_12998 = 6'h12 == _T_10211_40; // @[Mux.scala 46:19:@11032.4]
  assign _T_12999 = _T_12998 ? _T_9260_17 : _T_12997; // @[Mux.scala 46:16:@11033.4]
  assign _T_13000 = 6'h11 == _T_10211_40; // @[Mux.scala 46:19:@11034.4]
  assign _T_13001 = _T_13000 ? _T_9260_16 : _T_12999; // @[Mux.scala 46:16:@11035.4]
  assign _T_13002 = 6'h10 == _T_10211_40; // @[Mux.scala 46:19:@11036.4]
  assign _T_13003 = _T_13002 ? _T_9260_15 : _T_13001; // @[Mux.scala 46:16:@11037.4]
  assign _T_13004 = 6'hf == _T_10211_40; // @[Mux.scala 46:19:@11038.4]
  assign _T_13005 = _T_13004 ? _T_9260_14 : _T_13003; // @[Mux.scala 46:16:@11039.4]
  assign _T_13006 = 6'he == _T_10211_40; // @[Mux.scala 46:19:@11040.4]
  assign _T_13007 = _T_13006 ? _T_9260_13 : _T_13005; // @[Mux.scala 46:16:@11041.4]
  assign _T_13008 = 6'hd == _T_10211_40; // @[Mux.scala 46:19:@11042.4]
  assign _T_13009 = _T_13008 ? _T_9260_12 : _T_13007; // @[Mux.scala 46:16:@11043.4]
  assign _T_13010 = 6'hc == _T_10211_40; // @[Mux.scala 46:19:@11044.4]
  assign _T_13011 = _T_13010 ? _T_9260_11 : _T_13009; // @[Mux.scala 46:16:@11045.4]
  assign _T_13012 = 6'hb == _T_10211_40; // @[Mux.scala 46:19:@11046.4]
  assign _T_13013 = _T_13012 ? _T_9260_10 : _T_13011; // @[Mux.scala 46:16:@11047.4]
  assign _T_13014 = 6'ha == _T_10211_40; // @[Mux.scala 46:19:@11048.4]
  assign _T_13015 = _T_13014 ? _T_9260_9 : _T_13013; // @[Mux.scala 46:16:@11049.4]
  assign _T_13016 = 6'h9 == _T_10211_40; // @[Mux.scala 46:19:@11050.4]
  assign _T_13017 = _T_13016 ? _T_9260_8 : _T_13015; // @[Mux.scala 46:16:@11051.4]
  assign _T_13018 = 6'h8 == _T_10211_40; // @[Mux.scala 46:19:@11052.4]
  assign _T_13019 = _T_13018 ? _T_9260_7 : _T_13017; // @[Mux.scala 46:16:@11053.4]
  assign _T_13020 = 6'h7 == _T_10211_40; // @[Mux.scala 46:19:@11054.4]
  assign _T_13021 = _T_13020 ? _T_9260_6 : _T_13019; // @[Mux.scala 46:16:@11055.4]
  assign _T_13022 = 6'h6 == _T_10211_40; // @[Mux.scala 46:19:@11056.4]
  assign _T_13023 = _T_13022 ? _T_9260_5 : _T_13021; // @[Mux.scala 46:16:@11057.4]
  assign _T_13024 = 6'h5 == _T_10211_40; // @[Mux.scala 46:19:@11058.4]
  assign _T_13025 = _T_13024 ? _T_9260_4 : _T_13023; // @[Mux.scala 46:16:@11059.4]
  assign _T_13026 = 6'h4 == _T_10211_40; // @[Mux.scala 46:19:@11060.4]
  assign _T_13027 = _T_13026 ? _T_9260_3 : _T_13025; // @[Mux.scala 46:16:@11061.4]
  assign _T_13028 = 6'h3 == _T_10211_40; // @[Mux.scala 46:19:@11062.4]
  assign _T_13029 = _T_13028 ? _T_9260_2 : _T_13027; // @[Mux.scala 46:16:@11063.4]
  assign _T_13030 = 6'h2 == _T_10211_40; // @[Mux.scala 46:19:@11064.4]
  assign _T_13031 = _T_13030 ? _T_9260_1 : _T_13029; // @[Mux.scala 46:16:@11065.4]
  assign _T_13032 = 6'h1 == _T_10211_40; // @[Mux.scala 46:19:@11066.4]
  assign _T_13033 = _T_13032 ? _T_9260_0 : _T_13031; // @[Mux.scala 46:16:@11067.4]
  assign _T_13077 = 6'h2a == _T_10211_41; // @[Mux.scala 46:19:@11069.4]
  assign _T_13078 = _T_13077 ? _T_9260_41 : 8'h0; // @[Mux.scala 46:16:@11070.4]
  assign _T_13079 = 6'h29 == _T_10211_41; // @[Mux.scala 46:19:@11071.4]
  assign _T_13080 = _T_13079 ? _T_9260_40 : _T_13078; // @[Mux.scala 46:16:@11072.4]
  assign _T_13081 = 6'h28 == _T_10211_41; // @[Mux.scala 46:19:@11073.4]
  assign _T_13082 = _T_13081 ? _T_9260_39 : _T_13080; // @[Mux.scala 46:16:@11074.4]
  assign _T_13083 = 6'h27 == _T_10211_41; // @[Mux.scala 46:19:@11075.4]
  assign _T_13084 = _T_13083 ? _T_9260_38 : _T_13082; // @[Mux.scala 46:16:@11076.4]
  assign _T_13085 = 6'h26 == _T_10211_41; // @[Mux.scala 46:19:@11077.4]
  assign _T_13086 = _T_13085 ? _T_9260_37 : _T_13084; // @[Mux.scala 46:16:@11078.4]
  assign _T_13087 = 6'h25 == _T_10211_41; // @[Mux.scala 46:19:@11079.4]
  assign _T_13088 = _T_13087 ? _T_9260_36 : _T_13086; // @[Mux.scala 46:16:@11080.4]
  assign _T_13089 = 6'h24 == _T_10211_41; // @[Mux.scala 46:19:@11081.4]
  assign _T_13090 = _T_13089 ? _T_9260_35 : _T_13088; // @[Mux.scala 46:16:@11082.4]
  assign _T_13091 = 6'h23 == _T_10211_41; // @[Mux.scala 46:19:@11083.4]
  assign _T_13092 = _T_13091 ? _T_9260_34 : _T_13090; // @[Mux.scala 46:16:@11084.4]
  assign _T_13093 = 6'h22 == _T_10211_41; // @[Mux.scala 46:19:@11085.4]
  assign _T_13094 = _T_13093 ? _T_9260_33 : _T_13092; // @[Mux.scala 46:16:@11086.4]
  assign _T_13095 = 6'h21 == _T_10211_41; // @[Mux.scala 46:19:@11087.4]
  assign _T_13096 = _T_13095 ? _T_9260_32 : _T_13094; // @[Mux.scala 46:16:@11088.4]
  assign _T_13097 = 6'h20 == _T_10211_41; // @[Mux.scala 46:19:@11089.4]
  assign _T_13098 = _T_13097 ? _T_9260_31 : _T_13096; // @[Mux.scala 46:16:@11090.4]
  assign _T_13099 = 6'h1f == _T_10211_41; // @[Mux.scala 46:19:@11091.4]
  assign _T_13100 = _T_13099 ? _T_9260_30 : _T_13098; // @[Mux.scala 46:16:@11092.4]
  assign _T_13101 = 6'h1e == _T_10211_41; // @[Mux.scala 46:19:@11093.4]
  assign _T_13102 = _T_13101 ? _T_9260_29 : _T_13100; // @[Mux.scala 46:16:@11094.4]
  assign _T_13103 = 6'h1d == _T_10211_41; // @[Mux.scala 46:19:@11095.4]
  assign _T_13104 = _T_13103 ? _T_9260_28 : _T_13102; // @[Mux.scala 46:16:@11096.4]
  assign _T_13105 = 6'h1c == _T_10211_41; // @[Mux.scala 46:19:@11097.4]
  assign _T_13106 = _T_13105 ? _T_9260_27 : _T_13104; // @[Mux.scala 46:16:@11098.4]
  assign _T_13107 = 6'h1b == _T_10211_41; // @[Mux.scala 46:19:@11099.4]
  assign _T_13108 = _T_13107 ? _T_9260_26 : _T_13106; // @[Mux.scala 46:16:@11100.4]
  assign _T_13109 = 6'h1a == _T_10211_41; // @[Mux.scala 46:19:@11101.4]
  assign _T_13110 = _T_13109 ? _T_9260_25 : _T_13108; // @[Mux.scala 46:16:@11102.4]
  assign _T_13111 = 6'h19 == _T_10211_41; // @[Mux.scala 46:19:@11103.4]
  assign _T_13112 = _T_13111 ? _T_9260_24 : _T_13110; // @[Mux.scala 46:16:@11104.4]
  assign _T_13113 = 6'h18 == _T_10211_41; // @[Mux.scala 46:19:@11105.4]
  assign _T_13114 = _T_13113 ? _T_9260_23 : _T_13112; // @[Mux.scala 46:16:@11106.4]
  assign _T_13115 = 6'h17 == _T_10211_41; // @[Mux.scala 46:19:@11107.4]
  assign _T_13116 = _T_13115 ? _T_9260_22 : _T_13114; // @[Mux.scala 46:16:@11108.4]
  assign _T_13117 = 6'h16 == _T_10211_41; // @[Mux.scala 46:19:@11109.4]
  assign _T_13118 = _T_13117 ? _T_9260_21 : _T_13116; // @[Mux.scala 46:16:@11110.4]
  assign _T_13119 = 6'h15 == _T_10211_41; // @[Mux.scala 46:19:@11111.4]
  assign _T_13120 = _T_13119 ? _T_9260_20 : _T_13118; // @[Mux.scala 46:16:@11112.4]
  assign _T_13121 = 6'h14 == _T_10211_41; // @[Mux.scala 46:19:@11113.4]
  assign _T_13122 = _T_13121 ? _T_9260_19 : _T_13120; // @[Mux.scala 46:16:@11114.4]
  assign _T_13123 = 6'h13 == _T_10211_41; // @[Mux.scala 46:19:@11115.4]
  assign _T_13124 = _T_13123 ? _T_9260_18 : _T_13122; // @[Mux.scala 46:16:@11116.4]
  assign _T_13125 = 6'h12 == _T_10211_41; // @[Mux.scala 46:19:@11117.4]
  assign _T_13126 = _T_13125 ? _T_9260_17 : _T_13124; // @[Mux.scala 46:16:@11118.4]
  assign _T_13127 = 6'h11 == _T_10211_41; // @[Mux.scala 46:19:@11119.4]
  assign _T_13128 = _T_13127 ? _T_9260_16 : _T_13126; // @[Mux.scala 46:16:@11120.4]
  assign _T_13129 = 6'h10 == _T_10211_41; // @[Mux.scala 46:19:@11121.4]
  assign _T_13130 = _T_13129 ? _T_9260_15 : _T_13128; // @[Mux.scala 46:16:@11122.4]
  assign _T_13131 = 6'hf == _T_10211_41; // @[Mux.scala 46:19:@11123.4]
  assign _T_13132 = _T_13131 ? _T_9260_14 : _T_13130; // @[Mux.scala 46:16:@11124.4]
  assign _T_13133 = 6'he == _T_10211_41; // @[Mux.scala 46:19:@11125.4]
  assign _T_13134 = _T_13133 ? _T_9260_13 : _T_13132; // @[Mux.scala 46:16:@11126.4]
  assign _T_13135 = 6'hd == _T_10211_41; // @[Mux.scala 46:19:@11127.4]
  assign _T_13136 = _T_13135 ? _T_9260_12 : _T_13134; // @[Mux.scala 46:16:@11128.4]
  assign _T_13137 = 6'hc == _T_10211_41; // @[Mux.scala 46:19:@11129.4]
  assign _T_13138 = _T_13137 ? _T_9260_11 : _T_13136; // @[Mux.scala 46:16:@11130.4]
  assign _T_13139 = 6'hb == _T_10211_41; // @[Mux.scala 46:19:@11131.4]
  assign _T_13140 = _T_13139 ? _T_9260_10 : _T_13138; // @[Mux.scala 46:16:@11132.4]
  assign _T_13141 = 6'ha == _T_10211_41; // @[Mux.scala 46:19:@11133.4]
  assign _T_13142 = _T_13141 ? _T_9260_9 : _T_13140; // @[Mux.scala 46:16:@11134.4]
  assign _T_13143 = 6'h9 == _T_10211_41; // @[Mux.scala 46:19:@11135.4]
  assign _T_13144 = _T_13143 ? _T_9260_8 : _T_13142; // @[Mux.scala 46:16:@11136.4]
  assign _T_13145 = 6'h8 == _T_10211_41; // @[Mux.scala 46:19:@11137.4]
  assign _T_13146 = _T_13145 ? _T_9260_7 : _T_13144; // @[Mux.scala 46:16:@11138.4]
  assign _T_13147 = 6'h7 == _T_10211_41; // @[Mux.scala 46:19:@11139.4]
  assign _T_13148 = _T_13147 ? _T_9260_6 : _T_13146; // @[Mux.scala 46:16:@11140.4]
  assign _T_13149 = 6'h6 == _T_10211_41; // @[Mux.scala 46:19:@11141.4]
  assign _T_13150 = _T_13149 ? _T_9260_5 : _T_13148; // @[Mux.scala 46:16:@11142.4]
  assign _T_13151 = 6'h5 == _T_10211_41; // @[Mux.scala 46:19:@11143.4]
  assign _T_13152 = _T_13151 ? _T_9260_4 : _T_13150; // @[Mux.scala 46:16:@11144.4]
  assign _T_13153 = 6'h4 == _T_10211_41; // @[Mux.scala 46:19:@11145.4]
  assign _T_13154 = _T_13153 ? _T_9260_3 : _T_13152; // @[Mux.scala 46:16:@11146.4]
  assign _T_13155 = 6'h3 == _T_10211_41; // @[Mux.scala 46:19:@11147.4]
  assign _T_13156 = _T_13155 ? _T_9260_2 : _T_13154; // @[Mux.scala 46:16:@11148.4]
  assign _T_13157 = 6'h2 == _T_10211_41; // @[Mux.scala 46:19:@11149.4]
  assign _T_13158 = _T_13157 ? _T_9260_1 : _T_13156; // @[Mux.scala 46:16:@11150.4]
  assign _T_13159 = 6'h1 == _T_10211_41; // @[Mux.scala 46:19:@11151.4]
  assign _T_13160 = _T_13159 ? _T_9260_0 : _T_13158; // @[Mux.scala 46:16:@11152.4]
  assign _T_13205 = 6'h2b == _T_10211_42; // @[Mux.scala 46:19:@11154.4]
  assign _T_13206 = _T_13205 ? _T_9260_42 : 8'h0; // @[Mux.scala 46:16:@11155.4]
  assign _T_13207 = 6'h2a == _T_10211_42; // @[Mux.scala 46:19:@11156.4]
  assign _T_13208 = _T_13207 ? _T_9260_41 : _T_13206; // @[Mux.scala 46:16:@11157.4]
  assign _T_13209 = 6'h29 == _T_10211_42; // @[Mux.scala 46:19:@11158.4]
  assign _T_13210 = _T_13209 ? _T_9260_40 : _T_13208; // @[Mux.scala 46:16:@11159.4]
  assign _T_13211 = 6'h28 == _T_10211_42; // @[Mux.scala 46:19:@11160.4]
  assign _T_13212 = _T_13211 ? _T_9260_39 : _T_13210; // @[Mux.scala 46:16:@11161.4]
  assign _T_13213 = 6'h27 == _T_10211_42; // @[Mux.scala 46:19:@11162.4]
  assign _T_13214 = _T_13213 ? _T_9260_38 : _T_13212; // @[Mux.scala 46:16:@11163.4]
  assign _T_13215 = 6'h26 == _T_10211_42; // @[Mux.scala 46:19:@11164.4]
  assign _T_13216 = _T_13215 ? _T_9260_37 : _T_13214; // @[Mux.scala 46:16:@11165.4]
  assign _T_13217 = 6'h25 == _T_10211_42; // @[Mux.scala 46:19:@11166.4]
  assign _T_13218 = _T_13217 ? _T_9260_36 : _T_13216; // @[Mux.scala 46:16:@11167.4]
  assign _T_13219 = 6'h24 == _T_10211_42; // @[Mux.scala 46:19:@11168.4]
  assign _T_13220 = _T_13219 ? _T_9260_35 : _T_13218; // @[Mux.scala 46:16:@11169.4]
  assign _T_13221 = 6'h23 == _T_10211_42; // @[Mux.scala 46:19:@11170.4]
  assign _T_13222 = _T_13221 ? _T_9260_34 : _T_13220; // @[Mux.scala 46:16:@11171.4]
  assign _T_13223 = 6'h22 == _T_10211_42; // @[Mux.scala 46:19:@11172.4]
  assign _T_13224 = _T_13223 ? _T_9260_33 : _T_13222; // @[Mux.scala 46:16:@11173.4]
  assign _T_13225 = 6'h21 == _T_10211_42; // @[Mux.scala 46:19:@11174.4]
  assign _T_13226 = _T_13225 ? _T_9260_32 : _T_13224; // @[Mux.scala 46:16:@11175.4]
  assign _T_13227 = 6'h20 == _T_10211_42; // @[Mux.scala 46:19:@11176.4]
  assign _T_13228 = _T_13227 ? _T_9260_31 : _T_13226; // @[Mux.scala 46:16:@11177.4]
  assign _T_13229 = 6'h1f == _T_10211_42; // @[Mux.scala 46:19:@11178.4]
  assign _T_13230 = _T_13229 ? _T_9260_30 : _T_13228; // @[Mux.scala 46:16:@11179.4]
  assign _T_13231 = 6'h1e == _T_10211_42; // @[Mux.scala 46:19:@11180.4]
  assign _T_13232 = _T_13231 ? _T_9260_29 : _T_13230; // @[Mux.scala 46:16:@11181.4]
  assign _T_13233 = 6'h1d == _T_10211_42; // @[Mux.scala 46:19:@11182.4]
  assign _T_13234 = _T_13233 ? _T_9260_28 : _T_13232; // @[Mux.scala 46:16:@11183.4]
  assign _T_13235 = 6'h1c == _T_10211_42; // @[Mux.scala 46:19:@11184.4]
  assign _T_13236 = _T_13235 ? _T_9260_27 : _T_13234; // @[Mux.scala 46:16:@11185.4]
  assign _T_13237 = 6'h1b == _T_10211_42; // @[Mux.scala 46:19:@11186.4]
  assign _T_13238 = _T_13237 ? _T_9260_26 : _T_13236; // @[Mux.scala 46:16:@11187.4]
  assign _T_13239 = 6'h1a == _T_10211_42; // @[Mux.scala 46:19:@11188.4]
  assign _T_13240 = _T_13239 ? _T_9260_25 : _T_13238; // @[Mux.scala 46:16:@11189.4]
  assign _T_13241 = 6'h19 == _T_10211_42; // @[Mux.scala 46:19:@11190.4]
  assign _T_13242 = _T_13241 ? _T_9260_24 : _T_13240; // @[Mux.scala 46:16:@11191.4]
  assign _T_13243 = 6'h18 == _T_10211_42; // @[Mux.scala 46:19:@11192.4]
  assign _T_13244 = _T_13243 ? _T_9260_23 : _T_13242; // @[Mux.scala 46:16:@11193.4]
  assign _T_13245 = 6'h17 == _T_10211_42; // @[Mux.scala 46:19:@11194.4]
  assign _T_13246 = _T_13245 ? _T_9260_22 : _T_13244; // @[Mux.scala 46:16:@11195.4]
  assign _T_13247 = 6'h16 == _T_10211_42; // @[Mux.scala 46:19:@11196.4]
  assign _T_13248 = _T_13247 ? _T_9260_21 : _T_13246; // @[Mux.scala 46:16:@11197.4]
  assign _T_13249 = 6'h15 == _T_10211_42; // @[Mux.scala 46:19:@11198.4]
  assign _T_13250 = _T_13249 ? _T_9260_20 : _T_13248; // @[Mux.scala 46:16:@11199.4]
  assign _T_13251 = 6'h14 == _T_10211_42; // @[Mux.scala 46:19:@11200.4]
  assign _T_13252 = _T_13251 ? _T_9260_19 : _T_13250; // @[Mux.scala 46:16:@11201.4]
  assign _T_13253 = 6'h13 == _T_10211_42; // @[Mux.scala 46:19:@11202.4]
  assign _T_13254 = _T_13253 ? _T_9260_18 : _T_13252; // @[Mux.scala 46:16:@11203.4]
  assign _T_13255 = 6'h12 == _T_10211_42; // @[Mux.scala 46:19:@11204.4]
  assign _T_13256 = _T_13255 ? _T_9260_17 : _T_13254; // @[Mux.scala 46:16:@11205.4]
  assign _T_13257 = 6'h11 == _T_10211_42; // @[Mux.scala 46:19:@11206.4]
  assign _T_13258 = _T_13257 ? _T_9260_16 : _T_13256; // @[Mux.scala 46:16:@11207.4]
  assign _T_13259 = 6'h10 == _T_10211_42; // @[Mux.scala 46:19:@11208.4]
  assign _T_13260 = _T_13259 ? _T_9260_15 : _T_13258; // @[Mux.scala 46:16:@11209.4]
  assign _T_13261 = 6'hf == _T_10211_42; // @[Mux.scala 46:19:@11210.4]
  assign _T_13262 = _T_13261 ? _T_9260_14 : _T_13260; // @[Mux.scala 46:16:@11211.4]
  assign _T_13263 = 6'he == _T_10211_42; // @[Mux.scala 46:19:@11212.4]
  assign _T_13264 = _T_13263 ? _T_9260_13 : _T_13262; // @[Mux.scala 46:16:@11213.4]
  assign _T_13265 = 6'hd == _T_10211_42; // @[Mux.scala 46:19:@11214.4]
  assign _T_13266 = _T_13265 ? _T_9260_12 : _T_13264; // @[Mux.scala 46:16:@11215.4]
  assign _T_13267 = 6'hc == _T_10211_42; // @[Mux.scala 46:19:@11216.4]
  assign _T_13268 = _T_13267 ? _T_9260_11 : _T_13266; // @[Mux.scala 46:16:@11217.4]
  assign _T_13269 = 6'hb == _T_10211_42; // @[Mux.scala 46:19:@11218.4]
  assign _T_13270 = _T_13269 ? _T_9260_10 : _T_13268; // @[Mux.scala 46:16:@11219.4]
  assign _T_13271 = 6'ha == _T_10211_42; // @[Mux.scala 46:19:@11220.4]
  assign _T_13272 = _T_13271 ? _T_9260_9 : _T_13270; // @[Mux.scala 46:16:@11221.4]
  assign _T_13273 = 6'h9 == _T_10211_42; // @[Mux.scala 46:19:@11222.4]
  assign _T_13274 = _T_13273 ? _T_9260_8 : _T_13272; // @[Mux.scala 46:16:@11223.4]
  assign _T_13275 = 6'h8 == _T_10211_42; // @[Mux.scala 46:19:@11224.4]
  assign _T_13276 = _T_13275 ? _T_9260_7 : _T_13274; // @[Mux.scala 46:16:@11225.4]
  assign _T_13277 = 6'h7 == _T_10211_42; // @[Mux.scala 46:19:@11226.4]
  assign _T_13278 = _T_13277 ? _T_9260_6 : _T_13276; // @[Mux.scala 46:16:@11227.4]
  assign _T_13279 = 6'h6 == _T_10211_42; // @[Mux.scala 46:19:@11228.4]
  assign _T_13280 = _T_13279 ? _T_9260_5 : _T_13278; // @[Mux.scala 46:16:@11229.4]
  assign _T_13281 = 6'h5 == _T_10211_42; // @[Mux.scala 46:19:@11230.4]
  assign _T_13282 = _T_13281 ? _T_9260_4 : _T_13280; // @[Mux.scala 46:16:@11231.4]
  assign _T_13283 = 6'h4 == _T_10211_42; // @[Mux.scala 46:19:@11232.4]
  assign _T_13284 = _T_13283 ? _T_9260_3 : _T_13282; // @[Mux.scala 46:16:@11233.4]
  assign _T_13285 = 6'h3 == _T_10211_42; // @[Mux.scala 46:19:@11234.4]
  assign _T_13286 = _T_13285 ? _T_9260_2 : _T_13284; // @[Mux.scala 46:16:@11235.4]
  assign _T_13287 = 6'h2 == _T_10211_42; // @[Mux.scala 46:19:@11236.4]
  assign _T_13288 = _T_13287 ? _T_9260_1 : _T_13286; // @[Mux.scala 46:16:@11237.4]
  assign _T_13289 = 6'h1 == _T_10211_42; // @[Mux.scala 46:19:@11238.4]
  assign _T_13290 = _T_13289 ? _T_9260_0 : _T_13288; // @[Mux.scala 46:16:@11239.4]
  assign _T_13336 = 6'h2c == _T_10211_43; // @[Mux.scala 46:19:@11241.4]
  assign _T_13337 = _T_13336 ? _T_9260_43 : 8'h0; // @[Mux.scala 46:16:@11242.4]
  assign _T_13338 = 6'h2b == _T_10211_43; // @[Mux.scala 46:19:@11243.4]
  assign _T_13339 = _T_13338 ? _T_9260_42 : _T_13337; // @[Mux.scala 46:16:@11244.4]
  assign _T_13340 = 6'h2a == _T_10211_43; // @[Mux.scala 46:19:@11245.4]
  assign _T_13341 = _T_13340 ? _T_9260_41 : _T_13339; // @[Mux.scala 46:16:@11246.4]
  assign _T_13342 = 6'h29 == _T_10211_43; // @[Mux.scala 46:19:@11247.4]
  assign _T_13343 = _T_13342 ? _T_9260_40 : _T_13341; // @[Mux.scala 46:16:@11248.4]
  assign _T_13344 = 6'h28 == _T_10211_43; // @[Mux.scala 46:19:@11249.4]
  assign _T_13345 = _T_13344 ? _T_9260_39 : _T_13343; // @[Mux.scala 46:16:@11250.4]
  assign _T_13346 = 6'h27 == _T_10211_43; // @[Mux.scala 46:19:@11251.4]
  assign _T_13347 = _T_13346 ? _T_9260_38 : _T_13345; // @[Mux.scala 46:16:@11252.4]
  assign _T_13348 = 6'h26 == _T_10211_43; // @[Mux.scala 46:19:@11253.4]
  assign _T_13349 = _T_13348 ? _T_9260_37 : _T_13347; // @[Mux.scala 46:16:@11254.4]
  assign _T_13350 = 6'h25 == _T_10211_43; // @[Mux.scala 46:19:@11255.4]
  assign _T_13351 = _T_13350 ? _T_9260_36 : _T_13349; // @[Mux.scala 46:16:@11256.4]
  assign _T_13352 = 6'h24 == _T_10211_43; // @[Mux.scala 46:19:@11257.4]
  assign _T_13353 = _T_13352 ? _T_9260_35 : _T_13351; // @[Mux.scala 46:16:@11258.4]
  assign _T_13354 = 6'h23 == _T_10211_43; // @[Mux.scala 46:19:@11259.4]
  assign _T_13355 = _T_13354 ? _T_9260_34 : _T_13353; // @[Mux.scala 46:16:@11260.4]
  assign _T_13356 = 6'h22 == _T_10211_43; // @[Mux.scala 46:19:@11261.4]
  assign _T_13357 = _T_13356 ? _T_9260_33 : _T_13355; // @[Mux.scala 46:16:@11262.4]
  assign _T_13358 = 6'h21 == _T_10211_43; // @[Mux.scala 46:19:@11263.4]
  assign _T_13359 = _T_13358 ? _T_9260_32 : _T_13357; // @[Mux.scala 46:16:@11264.4]
  assign _T_13360 = 6'h20 == _T_10211_43; // @[Mux.scala 46:19:@11265.4]
  assign _T_13361 = _T_13360 ? _T_9260_31 : _T_13359; // @[Mux.scala 46:16:@11266.4]
  assign _T_13362 = 6'h1f == _T_10211_43; // @[Mux.scala 46:19:@11267.4]
  assign _T_13363 = _T_13362 ? _T_9260_30 : _T_13361; // @[Mux.scala 46:16:@11268.4]
  assign _T_13364 = 6'h1e == _T_10211_43; // @[Mux.scala 46:19:@11269.4]
  assign _T_13365 = _T_13364 ? _T_9260_29 : _T_13363; // @[Mux.scala 46:16:@11270.4]
  assign _T_13366 = 6'h1d == _T_10211_43; // @[Mux.scala 46:19:@11271.4]
  assign _T_13367 = _T_13366 ? _T_9260_28 : _T_13365; // @[Mux.scala 46:16:@11272.4]
  assign _T_13368 = 6'h1c == _T_10211_43; // @[Mux.scala 46:19:@11273.4]
  assign _T_13369 = _T_13368 ? _T_9260_27 : _T_13367; // @[Mux.scala 46:16:@11274.4]
  assign _T_13370 = 6'h1b == _T_10211_43; // @[Mux.scala 46:19:@11275.4]
  assign _T_13371 = _T_13370 ? _T_9260_26 : _T_13369; // @[Mux.scala 46:16:@11276.4]
  assign _T_13372 = 6'h1a == _T_10211_43; // @[Mux.scala 46:19:@11277.4]
  assign _T_13373 = _T_13372 ? _T_9260_25 : _T_13371; // @[Mux.scala 46:16:@11278.4]
  assign _T_13374 = 6'h19 == _T_10211_43; // @[Mux.scala 46:19:@11279.4]
  assign _T_13375 = _T_13374 ? _T_9260_24 : _T_13373; // @[Mux.scala 46:16:@11280.4]
  assign _T_13376 = 6'h18 == _T_10211_43; // @[Mux.scala 46:19:@11281.4]
  assign _T_13377 = _T_13376 ? _T_9260_23 : _T_13375; // @[Mux.scala 46:16:@11282.4]
  assign _T_13378 = 6'h17 == _T_10211_43; // @[Mux.scala 46:19:@11283.4]
  assign _T_13379 = _T_13378 ? _T_9260_22 : _T_13377; // @[Mux.scala 46:16:@11284.4]
  assign _T_13380 = 6'h16 == _T_10211_43; // @[Mux.scala 46:19:@11285.4]
  assign _T_13381 = _T_13380 ? _T_9260_21 : _T_13379; // @[Mux.scala 46:16:@11286.4]
  assign _T_13382 = 6'h15 == _T_10211_43; // @[Mux.scala 46:19:@11287.4]
  assign _T_13383 = _T_13382 ? _T_9260_20 : _T_13381; // @[Mux.scala 46:16:@11288.4]
  assign _T_13384 = 6'h14 == _T_10211_43; // @[Mux.scala 46:19:@11289.4]
  assign _T_13385 = _T_13384 ? _T_9260_19 : _T_13383; // @[Mux.scala 46:16:@11290.4]
  assign _T_13386 = 6'h13 == _T_10211_43; // @[Mux.scala 46:19:@11291.4]
  assign _T_13387 = _T_13386 ? _T_9260_18 : _T_13385; // @[Mux.scala 46:16:@11292.4]
  assign _T_13388 = 6'h12 == _T_10211_43; // @[Mux.scala 46:19:@11293.4]
  assign _T_13389 = _T_13388 ? _T_9260_17 : _T_13387; // @[Mux.scala 46:16:@11294.4]
  assign _T_13390 = 6'h11 == _T_10211_43; // @[Mux.scala 46:19:@11295.4]
  assign _T_13391 = _T_13390 ? _T_9260_16 : _T_13389; // @[Mux.scala 46:16:@11296.4]
  assign _T_13392 = 6'h10 == _T_10211_43; // @[Mux.scala 46:19:@11297.4]
  assign _T_13393 = _T_13392 ? _T_9260_15 : _T_13391; // @[Mux.scala 46:16:@11298.4]
  assign _T_13394 = 6'hf == _T_10211_43; // @[Mux.scala 46:19:@11299.4]
  assign _T_13395 = _T_13394 ? _T_9260_14 : _T_13393; // @[Mux.scala 46:16:@11300.4]
  assign _T_13396 = 6'he == _T_10211_43; // @[Mux.scala 46:19:@11301.4]
  assign _T_13397 = _T_13396 ? _T_9260_13 : _T_13395; // @[Mux.scala 46:16:@11302.4]
  assign _T_13398 = 6'hd == _T_10211_43; // @[Mux.scala 46:19:@11303.4]
  assign _T_13399 = _T_13398 ? _T_9260_12 : _T_13397; // @[Mux.scala 46:16:@11304.4]
  assign _T_13400 = 6'hc == _T_10211_43; // @[Mux.scala 46:19:@11305.4]
  assign _T_13401 = _T_13400 ? _T_9260_11 : _T_13399; // @[Mux.scala 46:16:@11306.4]
  assign _T_13402 = 6'hb == _T_10211_43; // @[Mux.scala 46:19:@11307.4]
  assign _T_13403 = _T_13402 ? _T_9260_10 : _T_13401; // @[Mux.scala 46:16:@11308.4]
  assign _T_13404 = 6'ha == _T_10211_43; // @[Mux.scala 46:19:@11309.4]
  assign _T_13405 = _T_13404 ? _T_9260_9 : _T_13403; // @[Mux.scala 46:16:@11310.4]
  assign _T_13406 = 6'h9 == _T_10211_43; // @[Mux.scala 46:19:@11311.4]
  assign _T_13407 = _T_13406 ? _T_9260_8 : _T_13405; // @[Mux.scala 46:16:@11312.4]
  assign _T_13408 = 6'h8 == _T_10211_43; // @[Mux.scala 46:19:@11313.4]
  assign _T_13409 = _T_13408 ? _T_9260_7 : _T_13407; // @[Mux.scala 46:16:@11314.4]
  assign _T_13410 = 6'h7 == _T_10211_43; // @[Mux.scala 46:19:@11315.4]
  assign _T_13411 = _T_13410 ? _T_9260_6 : _T_13409; // @[Mux.scala 46:16:@11316.4]
  assign _T_13412 = 6'h6 == _T_10211_43; // @[Mux.scala 46:19:@11317.4]
  assign _T_13413 = _T_13412 ? _T_9260_5 : _T_13411; // @[Mux.scala 46:16:@11318.4]
  assign _T_13414 = 6'h5 == _T_10211_43; // @[Mux.scala 46:19:@11319.4]
  assign _T_13415 = _T_13414 ? _T_9260_4 : _T_13413; // @[Mux.scala 46:16:@11320.4]
  assign _T_13416 = 6'h4 == _T_10211_43; // @[Mux.scala 46:19:@11321.4]
  assign _T_13417 = _T_13416 ? _T_9260_3 : _T_13415; // @[Mux.scala 46:16:@11322.4]
  assign _T_13418 = 6'h3 == _T_10211_43; // @[Mux.scala 46:19:@11323.4]
  assign _T_13419 = _T_13418 ? _T_9260_2 : _T_13417; // @[Mux.scala 46:16:@11324.4]
  assign _T_13420 = 6'h2 == _T_10211_43; // @[Mux.scala 46:19:@11325.4]
  assign _T_13421 = _T_13420 ? _T_9260_1 : _T_13419; // @[Mux.scala 46:16:@11326.4]
  assign _T_13422 = 6'h1 == _T_10211_43; // @[Mux.scala 46:19:@11327.4]
  assign _T_13423 = _T_13422 ? _T_9260_0 : _T_13421; // @[Mux.scala 46:16:@11328.4]
  assign _T_13470 = 6'h2d == _T_10211_44; // @[Mux.scala 46:19:@11330.4]
  assign _T_13471 = _T_13470 ? _T_9260_44 : 8'h0; // @[Mux.scala 46:16:@11331.4]
  assign _T_13472 = 6'h2c == _T_10211_44; // @[Mux.scala 46:19:@11332.4]
  assign _T_13473 = _T_13472 ? _T_9260_43 : _T_13471; // @[Mux.scala 46:16:@11333.4]
  assign _T_13474 = 6'h2b == _T_10211_44; // @[Mux.scala 46:19:@11334.4]
  assign _T_13475 = _T_13474 ? _T_9260_42 : _T_13473; // @[Mux.scala 46:16:@11335.4]
  assign _T_13476 = 6'h2a == _T_10211_44; // @[Mux.scala 46:19:@11336.4]
  assign _T_13477 = _T_13476 ? _T_9260_41 : _T_13475; // @[Mux.scala 46:16:@11337.4]
  assign _T_13478 = 6'h29 == _T_10211_44; // @[Mux.scala 46:19:@11338.4]
  assign _T_13479 = _T_13478 ? _T_9260_40 : _T_13477; // @[Mux.scala 46:16:@11339.4]
  assign _T_13480 = 6'h28 == _T_10211_44; // @[Mux.scala 46:19:@11340.4]
  assign _T_13481 = _T_13480 ? _T_9260_39 : _T_13479; // @[Mux.scala 46:16:@11341.4]
  assign _T_13482 = 6'h27 == _T_10211_44; // @[Mux.scala 46:19:@11342.4]
  assign _T_13483 = _T_13482 ? _T_9260_38 : _T_13481; // @[Mux.scala 46:16:@11343.4]
  assign _T_13484 = 6'h26 == _T_10211_44; // @[Mux.scala 46:19:@11344.4]
  assign _T_13485 = _T_13484 ? _T_9260_37 : _T_13483; // @[Mux.scala 46:16:@11345.4]
  assign _T_13486 = 6'h25 == _T_10211_44; // @[Mux.scala 46:19:@11346.4]
  assign _T_13487 = _T_13486 ? _T_9260_36 : _T_13485; // @[Mux.scala 46:16:@11347.4]
  assign _T_13488 = 6'h24 == _T_10211_44; // @[Mux.scala 46:19:@11348.4]
  assign _T_13489 = _T_13488 ? _T_9260_35 : _T_13487; // @[Mux.scala 46:16:@11349.4]
  assign _T_13490 = 6'h23 == _T_10211_44; // @[Mux.scala 46:19:@11350.4]
  assign _T_13491 = _T_13490 ? _T_9260_34 : _T_13489; // @[Mux.scala 46:16:@11351.4]
  assign _T_13492 = 6'h22 == _T_10211_44; // @[Mux.scala 46:19:@11352.4]
  assign _T_13493 = _T_13492 ? _T_9260_33 : _T_13491; // @[Mux.scala 46:16:@11353.4]
  assign _T_13494 = 6'h21 == _T_10211_44; // @[Mux.scala 46:19:@11354.4]
  assign _T_13495 = _T_13494 ? _T_9260_32 : _T_13493; // @[Mux.scala 46:16:@11355.4]
  assign _T_13496 = 6'h20 == _T_10211_44; // @[Mux.scala 46:19:@11356.4]
  assign _T_13497 = _T_13496 ? _T_9260_31 : _T_13495; // @[Mux.scala 46:16:@11357.4]
  assign _T_13498 = 6'h1f == _T_10211_44; // @[Mux.scala 46:19:@11358.4]
  assign _T_13499 = _T_13498 ? _T_9260_30 : _T_13497; // @[Mux.scala 46:16:@11359.4]
  assign _T_13500 = 6'h1e == _T_10211_44; // @[Mux.scala 46:19:@11360.4]
  assign _T_13501 = _T_13500 ? _T_9260_29 : _T_13499; // @[Mux.scala 46:16:@11361.4]
  assign _T_13502 = 6'h1d == _T_10211_44; // @[Mux.scala 46:19:@11362.4]
  assign _T_13503 = _T_13502 ? _T_9260_28 : _T_13501; // @[Mux.scala 46:16:@11363.4]
  assign _T_13504 = 6'h1c == _T_10211_44; // @[Mux.scala 46:19:@11364.4]
  assign _T_13505 = _T_13504 ? _T_9260_27 : _T_13503; // @[Mux.scala 46:16:@11365.4]
  assign _T_13506 = 6'h1b == _T_10211_44; // @[Mux.scala 46:19:@11366.4]
  assign _T_13507 = _T_13506 ? _T_9260_26 : _T_13505; // @[Mux.scala 46:16:@11367.4]
  assign _T_13508 = 6'h1a == _T_10211_44; // @[Mux.scala 46:19:@11368.4]
  assign _T_13509 = _T_13508 ? _T_9260_25 : _T_13507; // @[Mux.scala 46:16:@11369.4]
  assign _T_13510 = 6'h19 == _T_10211_44; // @[Mux.scala 46:19:@11370.4]
  assign _T_13511 = _T_13510 ? _T_9260_24 : _T_13509; // @[Mux.scala 46:16:@11371.4]
  assign _T_13512 = 6'h18 == _T_10211_44; // @[Mux.scala 46:19:@11372.4]
  assign _T_13513 = _T_13512 ? _T_9260_23 : _T_13511; // @[Mux.scala 46:16:@11373.4]
  assign _T_13514 = 6'h17 == _T_10211_44; // @[Mux.scala 46:19:@11374.4]
  assign _T_13515 = _T_13514 ? _T_9260_22 : _T_13513; // @[Mux.scala 46:16:@11375.4]
  assign _T_13516 = 6'h16 == _T_10211_44; // @[Mux.scala 46:19:@11376.4]
  assign _T_13517 = _T_13516 ? _T_9260_21 : _T_13515; // @[Mux.scala 46:16:@11377.4]
  assign _T_13518 = 6'h15 == _T_10211_44; // @[Mux.scala 46:19:@11378.4]
  assign _T_13519 = _T_13518 ? _T_9260_20 : _T_13517; // @[Mux.scala 46:16:@11379.4]
  assign _T_13520 = 6'h14 == _T_10211_44; // @[Mux.scala 46:19:@11380.4]
  assign _T_13521 = _T_13520 ? _T_9260_19 : _T_13519; // @[Mux.scala 46:16:@11381.4]
  assign _T_13522 = 6'h13 == _T_10211_44; // @[Mux.scala 46:19:@11382.4]
  assign _T_13523 = _T_13522 ? _T_9260_18 : _T_13521; // @[Mux.scala 46:16:@11383.4]
  assign _T_13524 = 6'h12 == _T_10211_44; // @[Mux.scala 46:19:@11384.4]
  assign _T_13525 = _T_13524 ? _T_9260_17 : _T_13523; // @[Mux.scala 46:16:@11385.4]
  assign _T_13526 = 6'h11 == _T_10211_44; // @[Mux.scala 46:19:@11386.4]
  assign _T_13527 = _T_13526 ? _T_9260_16 : _T_13525; // @[Mux.scala 46:16:@11387.4]
  assign _T_13528 = 6'h10 == _T_10211_44; // @[Mux.scala 46:19:@11388.4]
  assign _T_13529 = _T_13528 ? _T_9260_15 : _T_13527; // @[Mux.scala 46:16:@11389.4]
  assign _T_13530 = 6'hf == _T_10211_44; // @[Mux.scala 46:19:@11390.4]
  assign _T_13531 = _T_13530 ? _T_9260_14 : _T_13529; // @[Mux.scala 46:16:@11391.4]
  assign _T_13532 = 6'he == _T_10211_44; // @[Mux.scala 46:19:@11392.4]
  assign _T_13533 = _T_13532 ? _T_9260_13 : _T_13531; // @[Mux.scala 46:16:@11393.4]
  assign _T_13534 = 6'hd == _T_10211_44; // @[Mux.scala 46:19:@11394.4]
  assign _T_13535 = _T_13534 ? _T_9260_12 : _T_13533; // @[Mux.scala 46:16:@11395.4]
  assign _T_13536 = 6'hc == _T_10211_44; // @[Mux.scala 46:19:@11396.4]
  assign _T_13537 = _T_13536 ? _T_9260_11 : _T_13535; // @[Mux.scala 46:16:@11397.4]
  assign _T_13538 = 6'hb == _T_10211_44; // @[Mux.scala 46:19:@11398.4]
  assign _T_13539 = _T_13538 ? _T_9260_10 : _T_13537; // @[Mux.scala 46:16:@11399.4]
  assign _T_13540 = 6'ha == _T_10211_44; // @[Mux.scala 46:19:@11400.4]
  assign _T_13541 = _T_13540 ? _T_9260_9 : _T_13539; // @[Mux.scala 46:16:@11401.4]
  assign _T_13542 = 6'h9 == _T_10211_44; // @[Mux.scala 46:19:@11402.4]
  assign _T_13543 = _T_13542 ? _T_9260_8 : _T_13541; // @[Mux.scala 46:16:@11403.4]
  assign _T_13544 = 6'h8 == _T_10211_44; // @[Mux.scala 46:19:@11404.4]
  assign _T_13545 = _T_13544 ? _T_9260_7 : _T_13543; // @[Mux.scala 46:16:@11405.4]
  assign _T_13546 = 6'h7 == _T_10211_44; // @[Mux.scala 46:19:@11406.4]
  assign _T_13547 = _T_13546 ? _T_9260_6 : _T_13545; // @[Mux.scala 46:16:@11407.4]
  assign _T_13548 = 6'h6 == _T_10211_44; // @[Mux.scala 46:19:@11408.4]
  assign _T_13549 = _T_13548 ? _T_9260_5 : _T_13547; // @[Mux.scala 46:16:@11409.4]
  assign _T_13550 = 6'h5 == _T_10211_44; // @[Mux.scala 46:19:@11410.4]
  assign _T_13551 = _T_13550 ? _T_9260_4 : _T_13549; // @[Mux.scala 46:16:@11411.4]
  assign _T_13552 = 6'h4 == _T_10211_44; // @[Mux.scala 46:19:@11412.4]
  assign _T_13553 = _T_13552 ? _T_9260_3 : _T_13551; // @[Mux.scala 46:16:@11413.4]
  assign _T_13554 = 6'h3 == _T_10211_44; // @[Mux.scala 46:19:@11414.4]
  assign _T_13555 = _T_13554 ? _T_9260_2 : _T_13553; // @[Mux.scala 46:16:@11415.4]
  assign _T_13556 = 6'h2 == _T_10211_44; // @[Mux.scala 46:19:@11416.4]
  assign _T_13557 = _T_13556 ? _T_9260_1 : _T_13555; // @[Mux.scala 46:16:@11417.4]
  assign _T_13558 = 6'h1 == _T_10211_44; // @[Mux.scala 46:19:@11418.4]
  assign _T_13559 = _T_13558 ? _T_9260_0 : _T_13557; // @[Mux.scala 46:16:@11419.4]
  assign _T_13607 = 6'h2e == _T_10211_45; // @[Mux.scala 46:19:@11421.4]
  assign _T_13608 = _T_13607 ? _T_9260_45 : 8'h0; // @[Mux.scala 46:16:@11422.4]
  assign _T_13609 = 6'h2d == _T_10211_45; // @[Mux.scala 46:19:@11423.4]
  assign _T_13610 = _T_13609 ? _T_9260_44 : _T_13608; // @[Mux.scala 46:16:@11424.4]
  assign _T_13611 = 6'h2c == _T_10211_45; // @[Mux.scala 46:19:@11425.4]
  assign _T_13612 = _T_13611 ? _T_9260_43 : _T_13610; // @[Mux.scala 46:16:@11426.4]
  assign _T_13613 = 6'h2b == _T_10211_45; // @[Mux.scala 46:19:@11427.4]
  assign _T_13614 = _T_13613 ? _T_9260_42 : _T_13612; // @[Mux.scala 46:16:@11428.4]
  assign _T_13615 = 6'h2a == _T_10211_45; // @[Mux.scala 46:19:@11429.4]
  assign _T_13616 = _T_13615 ? _T_9260_41 : _T_13614; // @[Mux.scala 46:16:@11430.4]
  assign _T_13617 = 6'h29 == _T_10211_45; // @[Mux.scala 46:19:@11431.4]
  assign _T_13618 = _T_13617 ? _T_9260_40 : _T_13616; // @[Mux.scala 46:16:@11432.4]
  assign _T_13619 = 6'h28 == _T_10211_45; // @[Mux.scala 46:19:@11433.4]
  assign _T_13620 = _T_13619 ? _T_9260_39 : _T_13618; // @[Mux.scala 46:16:@11434.4]
  assign _T_13621 = 6'h27 == _T_10211_45; // @[Mux.scala 46:19:@11435.4]
  assign _T_13622 = _T_13621 ? _T_9260_38 : _T_13620; // @[Mux.scala 46:16:@11436.4]
  assign _T_13623 = 6'h26 == _T_10211_45; // @[Mux.scala 46:19:@11437.4]
  assign _T_13624 = _T_13623 ? _T_9260_37 : _T_13622; // @[Mux.scala 46:16:@11438.4]
  assign _T_13625 = 6'h25 == _T_10211_45; // @[Mux.scala 46:19:@11439.4]
  assign _T_13626 = _T_13625 ? _T_9260_36 : _T_13624; // @[Mux.scala 46:16:@11440.4]
  assign _T_13627 = 6'h24 == _T_10211_45; // @[Mux.scala 46:19:@11441.4]
  assign _T_13628 = _T_13627 ? _T_9260_35 : _T_13626; // @[Mux.scala 46:16:@11442.4]
  assign _T_13629 = 6'h23 == _T_10211_45; // @[Mux.scala 46:19:@11443.4]
  assign _T_13630 = _T_13629 ? _T_9260_34 : _T_13628; // @[Mux.scala 46:16:@11444.4]
  assign _T_13631 = 6'h22 == _T_10211_45; // @[Mux.scala 46:19:@11445.4]
  assign _T_13632 = _T_13631 ? _T_9260_33 : _T_13630; // @[Mux.scala 46:16:@11446.4]
  assign _T_13633 = 6'h21 == _T_10211_45; // @[Mux.scala 46:19:@11447.4]
  assign _T_13634 = _T_13633 ? _T_9260_32 : _T_13632; // @[Mux.scala 46:16:@11448.4]
  assign _T_13635 = 6'h20 == _T_10211_45; // @[Mux.scala 46:19:@11449.4]
  assign _T_13636 = _T_13635 ? _T_9260_31 : _T_13634; // @[Mux.scala 46:16:@11450.4]
  assign _T_13637 = 6'h1f == _T_10211_45; // @[Mux.scala 46:19:@11451.4]
  assign _T_13638 = _T_13637 ? _T_9260_30 : _T_13636; // @[Mux.scala 46:16:@11452.4]
  assign _T_13639 = 6'h1e == _T_10211_45; // @[Mux.scala 46:19:@11453.4]
  assign _T_13640 = _T_13639 ? _T_9260_29 : _T_13638; // @[Mux.scala 46:16:@11454.4]
  assign _T_13641 = 6'h1d == _T_10211_45; // @[Mux.scala 46:19:@11455.4]
  assign _T_13642 = _T_13641 ? _T_9260_28 : _T_13640; // @[Mux.scala 46:16:@11456.4]
  assign _T_13643 = 6'h1c == _T_10211_45; // @[Mux.scala 46:19:@11457.4]
  assign _T_13644 = _T_13643 ? _T_9260_27 : _T_13642; // @[Mux.scala 46:16:@11458.4]
  assign _T_13645 = 6'h1b == _T_10211_45; // @[Mux.scala 46:19:@11459.4]
  assign _T_13646 = _T_13645 ? _T_9260_26 : _T_13644; // @[Mux.scala 46:16:@11460.4]
  assign _T_13647 = 6'h1a == _T_10211_45; // @[Mux.scala 46:19:@11461.4]
  assign _T_13648 = _T_13647 ? _T_9260_25 : _T_13646; // @[Mux.scala 46:16:@11462.4]
  assign _T_13649 = 6'h19 == _T_10211_45; // @[Mux.scala 46:19:@11463.4]
  assign _T_13650 = _T_13649 ? _T_9260_24 : _T_13648; // @[Mux.scala 46:16:@11464.4]
  assign _T_13651 = 6'h18 == _T_10211_45; // @[Mux.scala 46:19:@11465.4]
  assign _T_13652 = _T_13651 ? _T_9260_23 : _T_13650; // @[Mux.scala 46:16:@11466.4]
  assign _T_13653 = 6'h17 == _T_10211_45; // @[Mux.scala 46:19:@11467.4]
  assign _T_13654 = _T_13653 ? _T_9260_22 : _T_13652; // @[Mux.scala 46:16:@11468.4]
  assign _T_13655 = 6'h16 == _T_10211_45; // @[Mux.scala 46:19:@11469.4]
  assign _T_13656 = _T_13655 ? _T_9260_21 : _T_13654; // @[Mux.scala 46:16:@11470.4]
  assign _T_13657 = 6'h15 == _T_10211_45; // @[Mux.scala 46:19:@11471.4]
  assign _T_13658 = _T_13657 ? _T_9260_20 : _T_13656; // @[Mux.scala 46:16:@11472.4]
  assign _T_13659 = 6'h14 == _T_10211_45; // @[Mux.scala 46:19:@11473.4]
  assign _T_13660 = _T_13659 ? _T_9260_19 : _T_13658; // @[Mux.scala 46:16:@11474.4]
  assign _T_13661 = 6'h13 == _T_10211_45; // @[Mux.scala 46:19:@11475.4]
  assign _T_13662 = _T_13661 ? _T_9260_18 : _T_13660; // @[Mux.scala 46:16:@11476.4]
  assign _T_13663 = 6'h12 == _T_10211_45; // @[Mux.scala 46:19:@11477.4]
  assign _T_13664 = _T_13663 ? _T_9260_17 : _T_13662; // @[Mux.scala 46:16:@11478.4]
  assign _T_13665 = 6'h11 == _T_10211_45; // @[Mux.scala 46:19:@11479.4]
  assign _T_13666 = _T_13665 ? _T_9260_16 : _T_13664; // @[Mux.scala 46:16:@11480.4]
  assign _T_13667 = 6'h10 == _T_10211_45; // @[Mux.scala 46:19:@11481.4]
  assign _T_13668 = _T_13667 ? _T_9260_15 : _T_13666; // @[Mux.scala 46:16:@11482.4]
  assign _T_13669 = 6'hf == _T_10211_45; // @[Mux.scala 46:19:@11483.4]
  assign _T_13670 = _T_13669 ? _T_9260_14 : _T_13668; // @[Mux.scala 46:16:@11484.4]
  assign _T_13671 = 6'he == _T_10211_45; // @[Mux.scala 46:19:@11485.4]
  assign _T_13672 = _T_13671 ? _T_9260_13 : _T_13670; // @[Mux.scala 46:16:@11486.4]
  assign _T_13673 = 6'hd == _T_10211_45; // @[Mux.scala 46:19:@11487.4]
  assign _T_13674 = _T_13673 ? _T_9260_12 : _T_13672; // @[Mux.scala 46:16:@11488.4]
  assign _T_13675 = 6'hc == _T_10211_45; // @[Mux.scala 46:19:@11489.4]
  assign _T_13676 = _T_13675 ? _T_9260_11 : _T_13674; // @[Mux.scala 46:16:@11490.4]
  assign _T_13677 = 6'hb == _T_10211_45; // @[Mux.scala 46:19:@11491.4]
  assign _T_13678 = _T_13677 ? _T_9260_10 : _T_13676; // @[Mux.scala 46:16:@11492.4]
  assign _T_13679 = 6'ha == _T_10211_45; // @[Mux.scala 46:19:@11493.4]
  assign _T_13680 = _T_13679 ? _T_9260_9 : _T_13678; // @[Mux.scala 46:16:@11494.4]
  assign _T_13681 = 6'h9 == _T_10211_45; // @[Mux.scala 46:19:@11495.4]
  assign _T_13682 = _T_13681 ? _T_9260_8 : _T_13680; // @[Mux.scala 46:16:@11496.4]
  assign _T_13683 = 6'h8 == _T_10211_45; // @[Mux.scala 46:19:@11497.4]
  assign _T_13684 = _T_13683 ? _T_9260_7 : _T_13682; // @[Mux.scala 46:16:@11498.4]
  assign _T_13685 = 6'h7 == _T_10211_45; // @[Mux.scala 46:19:@11499.4]
  assign _T_13686 = _T_13685 ? _T_9260_6 : _T_13684; // @[Mux.scala 46:16:@11500.4]
  assign _T_13687 = 6'h6 == _T_10211_45; // @[Mux.scala 46:19:@11501.4]
  assign _T_13688 = _T_13687 ? _T_9260_5 : _T_13686; // @[Mux.scala 46:16:@11502.4]
  assign _T_13689 = 6'h5 == _T_10211_45; // @[Mux.scala 46:19:@11503.4]
  assign _T_13690 = _T_13689 ? _T_9260_4 : _T_13688; // @[Mux.scala 46:16:@11504.4]
  assign _T_13691 = 6'h4 == _T_10211_45; // @[Mux.scala 46:19:@11505.4]
  assign _T_13692 = _T_13691 ? _T_9260_3 : _T_13690; // @[Mux.scala 46:16:@11506.4]
  assign _T_13693 = 6'h3 == _T_10211_45; // @[Mux.scala 46:19:@11507.4]
  assign _T_13694 = _T_13693 ? _T_9260_2 : _T_13692; // @[Mux.scala 46:16:@11508.4]
  assign _T_13695 = 6'h2 == _T_10211_45; // @[Mux.scala 46:19:@11509.4]
  assign _T_13696 = _T_13695 ? _T_9260_1 : _T_13694; // @[Mux.scala 46:16:@11510.4]
  assign _T_13697 = 6'h1 == _T_10211_45; // @[Mux.scala 46:19:@11511.4]
  assign _T_13698 = _T_13697 ? _T_9260_0 : _T_13696; // @[Mux.scala 46:16:@11512.4]
  assign _T_13747 = 6'h2f == _T_10211_46; // @[Mux.scala 46:19:@11514.4]
  assign _T_13748 = _T_13747 ? _T_9260_46 : 8'h0; // @[Mux.scala 46:16:@11515.4]
  assign _T_13749 = 6'h2e == _T_10211_46; // @[Mux.scala 46:19:@11516.4]
  assign _T_13750 = _T_13749 ? _T_9260_45 : _T_13748; // @[Mux.scala 46:16:@11517.4]
  assign _T_13751 = 6'h2d == _T_10211_46; // @[Mux.scala 46:19:@11518.4]
  assign _T_13752 = _T_13751 ? _T_9260_44 : _T_13750; // @[Mux.scala 46:16:@11519.4]
  assign _T_13753 = 6'h2c == _T_10211_46; // @[Mux.scala 46:19:@11520.4]
  assign _T_13754 = _T_13753 ? _T_9260_43 : _T_13752; // @[Mux.scala 46:16:@11521.4]
  assign _T_13755 = 6'h2b == _T_10211_46; // @[Mux.scala 46:19:@11522.4]
  assign _T_13756 = _T_13755 ? _T_9260_42 : _T_13754; // @[Mux.scala 46:16:@11523.4]
  assign _T_13757 = 6'h2a == _T_10211_46; // @[Mux.scala 46:19:@11524.4]
  assign _T_13758 = _T_13757 ? _T_9260_41 : _T_13756; // @[Mux.scala 46:16:@11525.4]
  assign _T_13759 = 6'h29 == _T_10211_46; // @[Mux.scala 46:19:@11526.4]
  assign _T_13760 = _T_13759 ? _T_9260_40 : _T_13758; // @[Mux.scala 46:16:@11527.4]
  assign _T_13761 = 6'h28 == _T_10211_46; // @[Mux.scala 46:19:@11528.4]
  assign _T_13762 = _T_13761 ? _T_9260_39 : _T_13760; // @[Mux.scala 46:16:@11529.4]
  assign _T_13763 = 6'h27 == _T_10211_46; // @[Mux.scala 46:19:@11530.4]
  assign _T_13764 = _T_13763 ? _T_9260_38 : _T_13762; // @[Mux.scala 46:16:@11531.4]
  assign _T_13765 = 6'h26 == _T_10211_46; // @[Mux.scala 46:19:@11532.4]
  assign _T_13766 = _T_13765 ? _T_9260_37 : _T_13764; // @[Mux.scala 46:16:@11533.4]
  assign _T_13767 = 6'h25 == _T_10211_46; // @[Mux.scala 46:19:@11534.4]
  assign _T_13768 = _T_13767 ? _T_9260_36 : _T_13766; // @[Mux.scala 46:16:@11535.4]
  assign _T_13769 = 6'h24 == _T_10211_46; // @[Mux.scala 46:19:@11536.4]
  assign _T_13770 = _T_13769 ? _T_9260_35 : _T_13768; // @[Mux.scala 46:16:@11537.4]
  assign _T_13771 = 6'h23 == _T_10211_46; // @[Mux.scala 46:19:@11538.4]
  assign _T_13772 = _T_13771 ? _T_9260_34 : _T_13770; // @[Mux.scala 46:16:@11539.4]
  assign _T_13773 = 6'h22 == _T_10211_46; // @[Mux.scala 46:19:@11540.4]
  assign _T_13774 = _T_13773 ? _T_9260_33 : _T_13772; // @[Mux.scala 46:16:@11541.4]
  assign _T_13775 = 6'h21 == _T_10211_46; // @[Mux.scala 46:19:@11542.4]
  assign _T_13776 = _T_13775 ? _T_9260_32 : _T_13774; // @[Mux.scala 46:16:@11543.4]
  assign _T_13777 = 6'h20 == _T_10211_46; // @[Mux.scala 46:19:@11544.4]
  assign _T_13778 = _T_13777 ? _T_9260_31 : _T_13776; // @[Mux.scala 46:16:@11545.4]
  assign _T_13779 = 6'h1f == _T_10211_46; // @[Mux.scala 46:19:@11546.4]
  assign _T_13780 = _T_13779 ? _T_9260_30 : _T_13778; // @[Mux.scala 46:16:@11547.4]
  assign _T_13781 = 6'h1e == _T_10211_46; // @[Mux.scala 46:19:@11548.4]
  assign _T_13782 = _T_13781 ? _T_9260_29 : _T_13780; // @[Mux.scala 46:16:@11549.4]
  assign _T_13783 = 6'h1d == _T_10211_46; // @[Mux.scala 46:19:@11550.4]
  assign _T_13784 = _T_13783 ? _T_9260_28 : _T_13782; // @[Mux.scala 46:16:@11551.4]
  assign _T_13785 = 6'h1c == _T_10211_46; // @[Mux.scala 46:19:@11552.4]
  assign _T_13786 = _T_13785 ? _T_9260_27 : _T_13784; // @[Mux.scala 46:16:@11553.4]
  assign _T_13787 = 6'h1b == _T_10211_46; // @[Mux.scala 46:19:@11554.4]
  assign _T_13788 = _T_13787 ? _T_9260_26 : _T_13786; // @[Mux.scala 46:16:@11555.4]
  assign _T_13789 = 6'h1a == _T_10211_46; // @[Mux.scala 46:19:@11556.4]
  assign _T_13790 = _T_13789 ? _T_9260_25 : _T_13788; // @[Mux.scala 46:16:@11557.4]
  assign _T_13791 = 6'h19 == _T_10211_46; // @[Mux.scala 46:19:@11558.4]
  assign _T_13792 = _T_13791 ? _T_9260_24 : _T_13790; // @[Mux.scala 46:16:@11559.4]
  assign _T_13793 = 6'h18 == _T_10211_46; // @[Mux.scala 46:19:@11560.4]
  assign _T_13794 = _T_13793 ? _T_9260_23 : _T_13792; // @[Mux.scala 46:16:@11561.4]
  assign _T_13795 = 6'h17 == _T_10211_46; // @[Mux.scala 46:19:@11562.4]
  assign _T_13796 = _T_13795 ? _T_9260_22 : _T_13794; // @[Mux.scala 46:16:@11563.4]
  assign _T_13797 = 6'h16 == _T_10211_46; // @[Mux.scala 46:19:@11564.4]
  assign _T_13798 = _T_13797 ? _T_9260_21 : _T_13796; // @[Mux.scala 46:16:@11565.4]
  assign _T_13799 = 6'h15 == _T_10211_46; // @[Mux.scala 46:19:@11566.4]
  assign _T_13800 = _T_13799 ? _T_9260_20 : _T_13798; // @[Mux.scala 46:16:@11567.4]
  assign _T_13801 = 6'h14 == _T_10211_46; // @[Mux.scala 46:19:@11568.4]
  assign _T_13802 = _T_13801 ? _T_9260_19 : _T_13800; // @[Mux.scala 46:16:@11569.4]
  assign _T_13803 = 6'h13 == _T_10211_46; // @[Mux.scala 46:19:@11570.4]
  assign _T_13804 = _T_13803 ? _T_9260_18 : _T_13802; // @[Mux.scala 46:16:@11571.4]
  assign _T_13805 = 6'h12 == _T_10211_46; // @[Mux.scala 46:19:@11572.4]
  assign _T_13806 = _T_13805 ? _T_9260_17 : _T_13804; // @[Mux.scala 46:16:@11573.4]
  assign _T_13807 = 6'h11 == _T_10211_46; // @[Mux.scala 46:19:@11574.4]
  assign _T_13808 = _T_13807 ? _T_9260_16 : _T_13806; // @[Mux.scala 46:16:@11575.4]
  assign _T_13809 = 6'h10 == _T_10211_46; // @[Mux.scala 46:19:@11576.4]
  assign _T_13810 = _T_13809 ? _T_9260_15 : _T_13808; // @[Mux.scala 46:16:@11577.4]
  assign _T_13811 = 6'hf == _T_10211_46; // @[Mux.scala 46:19:@11578.4]
  assign _T_13812 = _T_13811 ? _T_9260_14 : _T_13810; // @[Mux.scala 46:16:@11579.4]
  assign _T_13813 = 6'he == _T_10211_46; // @[Mux.scala 46:19:@11580.4]
  assign _T_13814 = _T_13813 ? _T_9260_13 : _T_13812; // @[Mux.scala 46:16:@11581.4]
  assign _T_13815 = 6'hd == _T_10211_46; // @[Mux.scala 46:19:@11582.4]
  assign _T_13816 = _T_13815 ? _T_9260_12 : _T_13814; // @[Mux.scala 46:16:@11583.4]
  assign _T_13817 = 6'hc == _T_10211_46; // @[Mux.scala 46:19:@11584.4]
  assign _T_13818 = _T_13817 ? _T_9260_11 : _T_13816; // @[Mux.scala 46:16:@11585.4]
  assign _T_13819 = 6'hb == _T_10211_46; // @[Mux.scala 46:19:@11586.4]
  assign _T_13820 = _T_13819 ? _T_9260_10 : _T_13818; // @[Mux.scala 46:16:@11587.4]
  assign _T_13821 = 6'ha == _T_10211_46; // @[Mux.scala 46:19:@11588.4]
  assign _T_13822 = _T_13821 ? _T_9260_9 : _T_13820; // @[Mux.scala 46:16:@11589.4]
  assign _T_13823 = 6'h9 == _T_10211_46; // @[Mux.scala 46:19:@11590.4]
  assign _T_13824 = _T_13823 ? _T_9260_8 : _T_13822; // @[Mux.scala 46:16:@11591.4]
  assign _T_13825 = 6'h8 == _T_10211_46; // @[Mux.scala 46:19:@11592.4]
  assign _T_13826 = _T_13825 ? _T_9260_7 : _T_13824; // @[Mux.scala 46:16:@11593.4]
  assign _T_13827 = 6'h7 == _T_10211_46; // @[Mux.scala 46:19:@11594.4]
  assign _T_13828 = _T_13827 ? _T_9260_6 : _T_13826; // @[Mux.scala 46:16:@11595.4]
  assign _T_13829 = 6'h6 == _T_10211_46; // @[Mux.scala 46:19:@11596.4]
  assign _T_13830 = _T_13829 ? _T_9260_5 : _T_13828; // @[Mux.scala 46:16:@11597.4]
  assign _T_13831 = 6'h5 == _T_10211_46; // @[Mux.scala 46:19:@11598.4]
  assign _T_13832 = _T_13831 ? _T_9260_4 : _T_13830; // @[Mux.scala 46:16:@11599.4]
  assign _T_13833 = 6'h4 == _T_10211_46; // @[Mux.scala 46:19:@11600.4]
  assign _T_13834 = _T_13833 ? _T_9260_3 : _T_13832; // @[Mux.scala 46:16:@11601.4]
  assign _T_13835 = 6'h3 == _T_10211_46; // @[Mux.scala 46:19:@11602.4]
  assign _T_13836 = _T_13835 ? _T_9260_2 : _T_13834; // @[Mux.scala 46:16:@11603.4]
  assign _T_13837 = 6'h2 == _T_10211_46; // @[Mux.scala 46:19:@11604.4]
  assign _T_13838 = _T_13837 ? _T_9260_1 : _T_13836; // @[Mux.scala 46:16:@11605.4]
  assign _T_13839 = 6'h1 == _T_10211_46; // @[Mux.scala 46:19:@11606.4]
  assign _T_13840 = _T_13839 ? _T_9260_0 : _T_13838; // @[Mux.scala 46:16:@11607.4]
  assign _T_13890 = 6'h30 == _T_10211_47; // @[Mux.scala 46:19:@11609.4]
  assign _T_13891 = _T_13890 ? _T_9260_47 : 8'h0; // @[Mux.scala 46:16:@11610.4]
  assign _T_13892 = 6'h2f == _T_10211_47; // @[Mux.scala 46:19:@11611.4]
  assign _T_13893 = _T_13892 ? _T_9260_46 : _T_13891; // @[Mux.scala 46:16:@11612.4]
  assign _T_13894 = 6'h2e == _T_10211_47; // @[Mux.scala 46:19:@11613.4]
  assign _T_13895 = _T_13894 ? _T_9260_45 : _T_13893; // @[Mux.scala 46:16:@11614.4]
  assign _T_13896 = 6'h2d == _T_10211_47; // @[Mux.scala 46:19:@11615.4]
  assign _T_13897 = _T_13896 ? _T_9260_44 : _T_13895; // @[Mux.scala 46:16:@11616.4]
  assign _T_13898 = 6'h2c == _T_10211_47; // @[Mux.scala 46:19:@11617.4]
  assign _T_13899 = _T_13898 ? _T_9260_43 : _T_13897; // @[Mux.scala 46:16:@11618.4]
  assign _T_13900 = 6'h2b == _T_10211_47; // @[Mux.scala 46:19:@11619.4]
  assign _T_13901 = _T_13900 ? _T_9260_42 : _T_13899; // @[Mux.scala 46:16:@11620.4]
  assign _T_13902 = 6'h2a == _T_10211_47; // @[Mux.scala 46:19:@11621.4]
  assign _T_13903 = _T_13902 ? _T_9260_41 : _T_13901; // @[Mux.scala 46:16:@11622.4]
  assign _T_13904 = 6'h29 == _T_10211_47; // @[Mux.scala 46:19:@11623.4]
  assign _T_13905 = _T_13904 ? _T_9260_40 : _T_13903; // @[Mux.scala 46:16:@11624.4]
  assign _T_13906 = 6'h28 == _T_10211_47; // @[Mux.scala 46:19:@11625.4]
  assign _T_13907 = _T_13906 ? _T_9260_39 : _T_13905; // @[Mux.scala 46:16:@11626.4]
  assign _T_13908 = 6'h27 == _T_10211_47; // @[Mux.scala 46:19:@11627.4]
  assign _T_13909 = _T_13908 ? _T_9260_38 : _T_13907; // @[Mux.scala 46:16:@11628.4]
  assign _T_13910 = 6'h26 == _T_10211_47; // @[Mux.scala 46:19:@11629.4]
  assign _T_13911 = _T_13910 ? _T_9260_37 : _T_13909; // @[Mux.scala 46:16:@11630.4]
  assign _T_13912 = 6'h25 == _T_10211_47; // @[Mux.scala 46:19:@11631.4]
  assign _T_13913 = _T_13912 ? _T_9260_36 : _T_13911; // @[Mux.scala 46:16:@11632.4]
  assign _T_13914 = 6'h24 == _T_10211_47; // @[Mux.scala 46:19:@11633.4]
  assign _T_13915 = _T_13914 ? _T_9260_35 : _T_13913; // @[Mux.scala 46:16:@11634.4]
  assign _T_13916 = 6'h23 == _T_10211_47; // @[Mux.scala 46:19:@11635.4]
  assign _T_13917 = _T_13916 ? _T_9260_34 : _T_13915; // @[Mux.scala 46:16:@11636.4]
  assign _T_13918 = 6'h22 == _T_10211_47; // @[Mux.scala 46:19:@11637.4]
  assign _T_13919 = _T_13918 ? _T_9260_33 : _T_13917; // @[Mux.scala 46:16:@11638.4]
  assign _T_13920 = 6'h21 == _T_10211_47; // @[Mux.scala 46:19:@11639.4]
  assign _T_13921 = _T_13920 ? _T_9260_32 : _T_13919; // @[Mux.scala 46:16:@11640.4]
  assign _T_13922 = 6'h20 == _T_10211_47; // @[Mux.scala 46:19:@11641.4]
  assign _T_13923 = _T_13922 ? _T_9260_31 : _T_13921; // @[Mux.scala 46:16:@11642.4]
  assign _T_13924 = 6'h1f == _T_10211_47; // @[Mux.scala 46:19:@11643.4]
  assign _T_13925 = _T_13924 ? _T_9260_30 : _T_13923; // @[Mux.scala 46:16:@11644.4]
  assign _T_13926 = 6'h1e == _T_10211_47; // @[Mux.scala 46:19:@11645.4]
  assign _T_13927 = _T_13926 ? _T_9260_29 : _T_13925; // @[Mux.scala 46:16:@11646.4]
  assign _T_13928 = 6'h1d == _T_10211_47; // @[Mux.scala 46:19:@11647.4]
  assign _T_13929 = _T_13928 ? _T_9260_28 : _T_13927; // @[Mux.scala 46:16:@11648.4]
  assign _T_13930 = 6'h1c == _T_10211_47; // @[Mux.scala 46:19:@11649.4]
  assign _T_13931 = _T_13930 ? _T_9260_27 : _T_13929; // @[Mux.scala 46:16:@11650.4]
  assign _T_13932 = 6'h1b == _T_10211_47; // @[Mux.scala 46:19:@11651.4]
  assign _T_13933 = _T_13932 ? _T_9260_26 : _T_13931; // @[Mux.scala 46:16:@11652.4]
  assign _T_13934 = 6'h1a == _T_10211_47; // @[Mux.scala 46:19:@11653.4]
  assign _T_13935 = _T_13934 ? _T_9260_25 : _T_13933; // @[Mux.scala 46:16:@11654.4]
  assign _T_13936 = 6'h19 == _T_10211_47; // @[Mux.scala 46:19:@11655.4]
  assign _T_13937 = _T_13936 ? _T_9260_24 : _T_13935; // @[Mux.scala 46:16:@11656.4]
  assign _T_13938 = 6'h18 == _T_10211_47; // @[Mux.scala 46:19:@11657.4]
  assign _T_13939 = _T_13938 ? _T_9260_23 : _T_13937; // @[Mux.scala 46:16:@11658.4]
  assign _T_13940 = 6'h17 == _T_10211_47; // @[Mux.scala 46:19:@11659.4]
  assign _T_13941 = _T_13940 ? _T_9260_22 : _T_13939; // @[Mux.scala 46:16:@11660.4]
  assign _T_13942 = 6'h16 == _T_10211_47; // @[Mux.scala 46:19:@11661.4]
  assign _T_13943 = _T_13942 ? _T_9260_21 : _T_13941; // @[Mux.scala 46:16:@11662.4]
  assign _T_13944 = 6'h15 == _T_10211_47; // @[Mux.scala 46:19:@11663.4]
  assign _T_13945 = _T_13944 ? _T_9260_20 : _T_13943; // @[Mux.scala 46:16:@11664.4]
  assign _T_13946 = 6'h14 == _T_10211_47; // @[Mux.scala 46:19:@11665.4]
  assign _T_13947 = _T_13946 ? _T_9260_19 : _T_13945; // @[Mux.scala 46:16:@11666.4]
  assign _T_13948 = 6'h13 == _T_10211_47; // @[Mux.scala 46:19:@11667.4]
  assign _T_13949 = _T_13948 ? _T_9260_18 : _T_13947; // @[Mux.scala 46:16:@11668.4]
  assign _T_13950 = 6'h12 == _T_10211_47; // @[Mux.scala 46:19:@11669.4]
  assign _T_13951 = _T_13950 ? _T_9260_17 : _T_13949; // @[Mux.scala 46:16:@11670.4]
  assign _T_13952 = 6'h11 == _T_10211_47; // @[Mux.scala 46:19:@11671.4]
  assign _T_13953 = _T_13952 ? _T_9260_16 : _T_13951; // @[Mux.scala 46:16:@11672.4]
  assign _T_13954 = 6'h10 == _T_10211_47; // @[Mux.scala 46:19:@11673.4]
  assign _T_13955 = _T_13954 ? _T_9260_15 : _T_13953; // @[Mux.scala 46:16:@11674.4]
  assign _T_13956 = 6'hf == _T_10211_47; // @[Mux.scala 46:19:@11675.4]
  assign _T_13957 = _T_13956 ? _T_9260_14 : _T_13955; // @[Mux.scala 46:16:@11676.4]
  assign _T_13958 = 6'he == _T_10211_47; // @[Mux.scala 46:19:@11677.4]
  assign _T_13959 = _T_13958 ? _T_9260_13 : _T_13957; // @[Mux.scala 46:16:@11678.4]
  assign _T_13960 = 6'hd == _T_10211_47; // @[Mux.scala 46:19:@11679.4]
  assign _T_13961 = _T_13960 ? _T_9260_12 : _T_13959; // @[Mux.scala 46:16:@11680.4]
  assign _T_13962 = 6'hc == _T_10211_47; // @[Mux.scala 46:19:@11681.4]
  assign _T_13963 = _T_13962 ? _T_9260_11 : _T_13961; // @[Mux.scala 46:16:@11682.4]
  assign _T_13964 = 6'hb == _T_10211_47; // @[Mux.scala 46:19:@11683.4]
  assign _T_13965 = _T_13964 ? _T_9260_10 : _T_13963; // @[Mux.scala 46:16:@11684.4]
  assign _T_13966 = 6'ha == _T_10211_47; // @[Mux.scala 46:19:@11685.4]
  assign _T_13967 = _T_13966 ? _T_9260_9 : _T_13965; // @[Mux.scala 46:16:@11686.4]
  assign _T_13968 = 6'h9 == _T_10211_47; // @[Mux.scala 46:19:@11687.4]
  assign _T_13969 = _T_13968 ? _T_9260_8 : _T_13967; // @[Mux.scala 46:16:@11688.4]
  assign _T_13970 = 6'h8 == _T_10211_47; // @[Mux.scala 46:19:@11689.4]
  assign _T_13971 = _T_13970 ? _T_9260_7 : _T_13969; // @[Mux.scala 46:16:@11690.4]
  assign _T_13972 = 6'h7 == _T_10211_47; // @[Mux.scala 46:19:@11691.4]
  assign _T_13973 = _T_13972 ? _T_9260_6 : _T_13971; // @[Mux.scala 46:16:@11692.4]
  assign _T_13974 = 6'h6 == _T_10211_47; // @[Mux.scala 46:19:@11693.4]
  assign _T_13975 = _T_13974 ? _T_9260_5 : _T_13973; // @[Mux.scala 46:16:@11694.4]
  assign _T_13976 = 6'h5 == _T_10211_47; // @[Mux.scala 46:19:@11695.4]
  assign _T_13977 = _T_13976 ? _T_9260_4 : _T_13975; // @[Mux.scala 46:16:@11696.4]
  assign _T_13978 = 6'h4 == _T_10211_47; // @[Mux.scala 46:19:@11697.4]
  assign _T_13979 = _T_13978 ? _T_9260_3 : _T_13977; // @[Mux.scala 46:16:@11698.4]
  assign _T_13980 = 6'h3 == _T_10211_47; // @[Mux.scala 46:19:@11699.4]
  assign _T_13981 = _T_13980 ? _T_9260_2 : _T_13979; // @[Mux.scala 46:16:@11700.4]
  assign _T_13982 = 6'h2 == _T_10211_47; // @[Mux.scala 46:19:@11701.4]
  assign _T_13983 = _T_13982 ? _T_9260_1 : _T_13981; // @[Mux.scala 46:16:@11702.4]
  assign _T_13984 = 6'h1 == _T_10211_47; // @[Mux.scala 46:19:@11703.4]
  assign _T_13985 = _T_13984 ? _T_9260_0 : _T_13983; // @[Mux.scala 46:16:@11704.4]
  assign _T_14036 = 6'h31 == _T_10211_48; // @[Mux.scala 46:19:@11706.4]
  assign _T_14037 = _T_14036 ? _T_9260_48 : 8'h0; // @[Mux.scala 46:16:@11707.4]
  assign _T_14038 = 6'h30 == _T_10211_48; // @[Mux.scala 46:19:@11708.4]
  assign _T_14039 = _T_14038 ? _T_9260_47 : _T_14037; // @[Mux.scala 46:16:@11709.4]
  assign _T_14040 = 6'h2f == _T_10211_48; // @[Mux.scala 46:19:@11710.4]
  assign _T_14041 = _T_14040 ? _T_9260_46 : _T_14039; // @[Mux.scala 46:16:@11711.4]
  assign _T_14042 = 6'h2e == _T_10211_48; // @[Mux.scala 46:19:@11712.4]
  assign _T_14043 = _T_14042 ? _T_9260_45 : _T_14041; // @[Mux.scala 46:16:@11713.4]
  assign _T_14044 = 6'h2d == _T_10211_48; // @[Mux.scala 46:19:@11714.4]
  assign _T_14045 = _T_14044 ? _T_9260_44 : _T_14043; // @[Mux.scala 46:16:@11715.4]
  assign _T_14046 = 6'h2c == _T_10211_48; // @[Mux.scala 46:19:@11716.4]
  assign _T_14047 = _T_14046 ? _T_9260_43 : _T_14045; // @[Mux.scala 46:16:@11717.4]
  assign _T_14048 = 6'h2b == _T_10211_48; // @[Mux.scala 46:19:@11718.4]
  assign _T_14049 = _T_14048 ? _T_9260_42 : _T_14047; // @[Mux.scala 46:16:@11719.4]
  assign _T_14050 = 6'h2a == _T_10211_48; // @[Mux.scala 46:19:@11720.4]
  assign _T_14051 = _T_14050 ? _T_9260_41 : _T_14049; // @[Mux.scala 46:16:@11721.4]
  assign _T_14052 = 6'h29 == _T_10211_48; // @[Mux.scala 46:19:@11722.4]
  assign _T_14053 = _T_14052 ? _T_9260_40 : _T_14051; // @[Mux.scala 46:16:@11723.4]
  assign _T_14054 = 6'h28 == _T_10211_48; // @[Mux.scala 46:19:@11724.4]
  assign _T_14055 = _T_14054 ? _T_9260_39 : _T_14053; // @[Mux.scala 46:16:@11725.4]
  assign _T_14056 = 6'h27 == _T_10211_48; // @[Mux.scala 46:19:@11726.4]
  assign _T_14057 = _T_14056 ? _T_9260_38 : _T_14055; // @[Mux.scala 46:16:@11727.4]
  assign _T_14058 = 6'h26 == _T_10211_48; // @[Mux.scala 46:19:@11728.4]
  assign _T_14059 = _T_14058 ? _T_9260_37 : _T_14057; // @[Mux.scala 46:16:@11729.4]
  assign _T_14060 = 6'h25 == _T_10211_48; // @[Mux.scala 46:19:@11730.4]
  assign _T_14061 = _T_14060 ? _T_9260_36 : _T_14059; // @[Mux.scala 46:16:@11731.4]
  assign _T_14062 = 6'h24 == _T_10211_48; // @[Mux.scala 46:19:@11732.4]
  assign _T_14063 = _T_14062 ? _T_9260_35 : _T_14061; // @[Mux.scala 46:16:@11733.4]
  assign _T_14064 = 6'h23 == _T_10211_48; // @[Mux.scala 46:19:@11734.4]
  assign _T_14065 = _T_14064 ? _T_9260_34 : _T_14063; // @[Mux.scala 46:16:@11735.4]
  assign _T_14066 = 6'h22 == _T_10211_48; // @[Mux.scala 46:19:@11736.4]
  assign _T_14067 = _T_14066 ? _T_9260_33 : _T_14065; // @[Mux.scala 46:16:@11737.4]
  assign _T_14068 = 6'h21 == _T_10211_48; // @[Mux.scala 46:19:@11738.4]
  assign _T_14069 = _T_14068 ? _T_9260_32 : _T_14067; // @[Mux.scala 46:16:@11739.4]
  assign _T_14070 = 6'h20 == _T_10211_48; // @[Mux.scala 46:19:@11740.4]
  assign _T_14071 = _T_14070 ? _T_9260_31 : _T_14069; // @[Mux.scala 46:16:@11741.4]
  assign _T_14072 = 6'h1f == _T_10211_48; // @[Mux.scala 46:19:@11742.4]
  assign _T_14073 = _T_14072 ? _T_9260_30 : _T_14071; // @[Mux.scala 46:16:@11743.4]
  assign _T_14074 = 6'h1e == _T_10211_48; // @[Mux.scala 46:19:@11744.4]
  assign _T_14075 = _T_14074 ? _T_9260_29 : _T_14073; // @[Mux.scala 46:16:@11745.4]
  assign _T_14076 = 6'h1d == _T_10211_48; // @[Mux.scala 46:19:@11746.4]
  assign _T_14077 = _T_14076 ? _T_9260_28 : _T_14075; // @[Mux.scala 46:16:@11747.4]
  assign _T_14078 = 6'h1c == _T_10211_48; // @[Mux.scala 46:19:@11748.4]
  assign _T_14079 = _T_14078 ? _T_9260_27 : _T_14077; // @[Mux.scala 46:16:@11749.4]
  assign _T_14080 = 6'h1b == _T_10211_48; // @[Mux.scala 46:19:@11750.4]
  assign _T_14081 = _T_14080 ? _T_9260_26 : _T_14079; // @[Mux.scala 46:16:@11751.4]
  assign _T_14082 = 6'h1a == _T_10211_48; // @[Mux.scala 46:19:@11752.4]
  assign _T_14083 = _T_14082 ? _T_9260_25 : _T_14081; // @[Mux.scala 46:16:@11753.4]
  assign _T_14084 = 6'h19 == _T_10211_48; // @[Mux.scala 46:19:@11754.4]
  assign _T_14085 = _T_14084 ? _T_9260_24 : _T_14083; // @[Mux.scala 46:16:@11755.4]
  assign _T_14086 = 6'h18 == _T_10211_48; // @[Mux.scala 46:19:@11756.4]
  assign _T_14087 = _T_14086 ? _T_9260_23 : _T_14085; // @[Mux.scala 46:16:@11757.4]
  assign _T_14088 = 6'h17 == _T_10211_48; // @[Mux.scala 46:19:@11758.4]
  assign _T_14089 = _T_14088 ? _T_9260_22 : _T_14087; // @[Mux.scala 46:16:@11759.4]
  assign _T_14090 = 6'h16 == _T_10211_48; // @[Mux.scala 46:19:@11760.4]
  assign _T_14091 = _T_14090 ? _T_9260_21 : _T_14089; // @[Mux.scala 46:16:@11761.4]
  assign _T_14092 = 6'h15 == _T_10211_48; // @[Mux.scala 46:19:@11762.4]
  assign _T_14093 = _T_14092 ? _T_9260_20 : _T_14091; // @[Mux.scala 46:16:@11763.4]
  assign _T_14094 = 6'h14 == _T_10211_48; // @[Mux.scala 46:19:@11764.4]
  assign _T_14095 = _T_14094 ? _T_9260_19 : _T_14093; // @[Mux.scala 46:16:@11765.4]
  assign _T_14096 = 6'h13 == _T_10211_48; // @[Mux.scala 46:19:@11766.4]
  assign _T_14097 = _T_14096 ? _T_9260_18 : _T_14095; // @[Mux.scala 46:16:@11767.4]
  assign _T_14098 = 6'h12 == _T_10211_48; // @[Mux.scala 46:19:@11768.4]
  assign _T_14099 = _T_14098 ? _T_9260_17 : _T_14097; // @[Mux.scala 46:16:@11769.4]
  assign _T_14100 = 6'h11 == _T_10211_48; // @[Mux.scala 46:19:@11770.4]
  assign _T_14101 = _T_14100 ? _T_9260_16 : _T_14099; // @[Mux.scala 46:16:@11771.4]
  assign _T_14102 = 6'h10 == _T_10211_48; // @[Mux.scala 46:19:@11772.4]
  assign _T_14103 = _T_14102 ? _T_9260_15 : _T_14101; // @[Mux.scala 46:16:@11773.4]
  assign _T_14104 = 6'hf == _T_10211_48; // @[Mux.scala 46:19:@11774.4]
  assign _T_14105 = _T_14104 ? _T_9260_14 : _T_14103; // @[Mux.scala 46:16:@11775.4]
  assign _T_14106 = 6'he == _T_10211_48; // @[Mux.scala 46:19:@11776.4]
  assign _T_14107 = _T_14106 ? _T_9260_13 : _T_14105; // @[Mux.scala 46:16:@11777.4]
  assign _T_14108 = 6'hd == _T_10211_48; // @[Mux.scala 46:19:@11778.4]
  assign _T_14109 = _T_14108 ? _T_9260_12 : _T_14107; // @[Mux.scala 46:16:@11779.4]
  assign _T_14110 = 6'hc == _T_10211_48; // @[Mux.scala 46:19:@11780.4]
  assign _T_14111 = _T_14110 ? _T_9260_11 : _T_14109; // @[Mux.scala 46:16:@11781.4]
  assign _T_14112 = 6'hb == _T_10211_48; // @[Mux.scala 46:19:@11782.4]
  assign _T_14113 = _T_14112 ? _T_9260_10 : _T_14111; // @[Mux.scala 46:16:@11783.4]
  assign _T_14114 = 6'ha == _T_10211_48; // @[Mux.scala 46:19:@11784.4]
  assign _T_14115 = _T_14114 ? _T_9260_9 : _T_14113; // @[Mux.scala 46:16:@11785.4]
  assign _T_14116 = 6'h9 == _T_10211_48; // @[Mux.scala 46:19:@11786.4]
  assign _T_14117 = _T_14116 ? _T_9260_8 : _T_14115; // @[Mux.scala 46:16:@11787.4]
  assign _T_14118 = 6'h8 == _T_10211_48; // @[Mux.scala 46:19:@11788.4]
  assign _T_14119 = _T_14118 ? _T_9260_7 : _T_14117; // @[Mux.scala 46:16:@11789.4]
  assign _T_14120 = 6'h7 == _T_10211_48; // @[Mux.scala 46:19:@11790.4]
  assign _T_14121 = _T_14120 ? _T_9260_6 : _T_14119; // @[Mux.scala 46:16:@11791.4]
  assign _T_14122 = 6'h6 == _T_10211_48; // @[Mux.scala 46:19:@11792.4]
  assign _T_14123 = _T_14122 ? _T_9260_5 : _T_14121; // @[Mux.scala 46:16:@11793.4]
  assign _T_14124 = 6'h5 == _T_10211_48; // @[Mux.scala 46:19:@11794.4]
  assign _T_14125 = _T_14124 ? _T_9260_4 : _T_14123; // @[Mux.scala 46:16:@11795.4]
  assign _T_14126 = 6'h4 == _T_10211_48; // @[Mux.scala 46:19:@11796.4]
  assign _T_14127 = _T_14126 ? _T_9260_3 : _T_14125; // @[Mux.scala 46:16:@11797.4]
  assign _T_14128 = 6'h3 == _T_10211_48; // @[Mux.scala 46:19:@11798.4]
  assign _T_14129 = _T_14128 ? _T_9260_2 : _T_14127; // @[Mux.scala 46:16:@11799.4]
  assign _T_14130 = 6'h2 == _T_10211_48; // @[Mux.scala 46:19:@11800.4]
  assign _T_14131 = _T_14130 ? _T_9260_1 : _T_14129; // @[Mux.scala 46:16:@11801.4]
  assign _T_14132 = 6'h1 == _T_10211_48; // @[Mux.scala 46:19:@11802.4]
  assign _T_14133 = _T_14132 ? _T_9260_0 : _T_14131; // @[Mux.scala 46:16:@11803.4]
  assign _T_14185 = 6'h32 == _T_10211_49; // @[Mux.scala 46:19:@11805.4]
  assign _T_14186 = _T_14185 ? _T_9260_49 : 8'h0; // @[Mux.scala 46:16:@11806.4]
  assign _T_14187 = 6'h31 == _T_10211_49; // @[Mux.scala 46:19:@11807.4]
  assign _T_14188 = _T_14187 ? _T_9260_48 : _T_14186; // @[Mux.scala 46:16:@11808.4]
  assign _T_14189 = 6'h30 == _T_10211_49; // @[Mux.scala 46:19:@11809.4]
  assign _T_14190 = _T_14189 ? _T_9260_47 : _T_14188; // @[Mux.scala 46:16:@11810.4]
  assign _T_14191 = 6'h2f == _T_10211_49; // @[Mux.scala 46:19:@11811.4]
  assign _T_14192 = _T_14191 ? _T_9260_46 : _T_14190; // @[Mux.scala 46:16:@11812.4]
  assign _T_14193 = 6'h2e == _T_10211_49; // @[Mux.scala 46:19:@11813.4]
  assign _T_14194 = _T_14193 ? _T_9260_45 : _T_14192; // @[Mux.scala 46:16:@11814.4]
  assign _T_14195 = 6'h2d == _T_10211_49; // @[Mux.scala 46:19:@11815.4]
  assign _T_14196 = _T_14195 ? _T_9260_44 : _T_14194; // @[Mux.scala 46:16:@11816.4]
  assign _T_14197 = 6'h2c == _T_10211_49; // @[Mux.scala 46:19:@11817.4]
  assign _T_14198 = _T_14197 ? _T_9260_43 : _T_14196; // @[Mux.scala 46:16:@11818.4]
  assign _T_14199 = 6'h2b == _T_10211_49; // @[Mux.scala 46:19:@11819.4]
  assign _T_14200 = _T_14199 ? _T_9260_42 : _T_14198; // @[Mux.scala 46:16:@11820.4]
  assign _T_14201 = 6'h2a == _T_10211_49; // @[Mux.scala 46:19:@11821.4]
  assign _T_14202 = _T_14201 ? _T_9260_41 : _T_14200; // @[Mux.scala 46:16:@11822.4]
  assign _T_14203 = 6'h29 == _T_10211_49; // @[Mux.scala 46:19:@11823.4]
  assign _T_14204 = _T_14203 ? _T_9260_40 : _T_14202; // @[Mux.scala 46:16:@11824.4]
  assign _T_14205 = 6'h28 == _T_10211_49; // @[Mux.scala 46:19:@11825.4]
  assign _T_14206 = _T_14205 ? _T_9260_39 : _T_14204; // @[Mux.scala 46:16:@11826.4]
  assign _T_14207 = 6'h27 == _T_10211_49; // @[Mux.scala 46:19:@11827.4]
  assign _T_14208 = _T_14207 ? _T_9260_38 : _T_14206; // @[Mux.scala 46:16:@11828.4]
  assign _T_14209 = 6'h26 == _T_10211_49; // @[Mux.scala 46:19:@11829.4]
  assign _T_14210 = _T_14209 ? _T_9260_37 : _T_14208; // @[Mux.scala 46:16:@11830.4]
  assign _T_14211 = 6'h25 == _T_10211_49; // @[Mux.scala 46:19:@11831.4]
  assign _T_14212 = _T_14211 ? _T_9260_36 : _T_14210; // @[Mux.scala 46:16:@11832.4]
  assign _T_14213 = 6'h24 == _T_10211_49; // @[Mux.scala 46:19:@11833.4]
  assign _T_14214 = _T_14213 ? _T_9260_35 : _T_14212; // @[Mux.scala 46:16:@11834.4]
  assign _T_14215 = 6'h23 == _T_10211_49; // @[Mux.scala 46:19:@11835.4]
  assign _T_14216 = _T_14215 ? _T_9260_34 : _T_14214; // @[Mux.scala 46:16:@11836.4]
  assign _T_14217 = 6'h22 == _T_10211_49; // @[Mux.scala 46:19:@11837.4]
  assign _T_14218 = _T_14217 ? _T_9260_33 : _T_14216; // @[Mux.scala 46:16:@11838.4]
  assign _T_14219 = 6'h21 == _T_10211_49; // @[Mux.scala 46:19:@11839.4]
  assign _T_14220 = _T_14219 ? _T_9260_32 : _T_14218; // @[Mux.scala 46:16:@11840.4]
  assign _T_14221 = 6'h20 == _T_10211_49; // @[Mux.scala 46:19:@11841.4]
  assign _T_14222 = _T_14221 ? _T_9260_31 : _T_14220; // @[Mux.scala 46:16:@11842.4]
  assign _T_14223 = 6'h1f == _T_10211_49; // @[Mux.scala 46:19:@11843.4]
  assign _T_14224 = _T_14223 ? _T_9260_30 : _T_14222; // @[Mux.scala 46:16:@11844.4]
  assign _T_14225 = 6'h1e == _T_10211_49; // @[Mux.scala 46:19:@11845.4]
  assign _T_14226 = _T_14225 ? _T_9260_29 : _T_14224; // @[Mux.scala 46:16:@11846.4]
  assign _T_14227 = 6'h1d == _T_10211_49; // @[Mux.scala 46:19:@11847.4]
  assign _T_14228 = _T_14227 ? _T_9260_28 : _T_14226; // @[Mux.scala 46:16:@11848.4]
  assign _T_14229 = 6'h1c == _T_10211_49; // @[Mux.scala 46:19:@11849.4]
  assign _T_14230 = _T_14229 ? _T_9260_27 : _T_14228; // @[Mux.scala 46:16:@11850.4]
  assign _T_14231 = 6'h1b == _T_10211_49; // @[Mux.scala 46:19:@11851.4]
  assign _T_14232 = _T_14231 ? _T_9260_26 : _T_14230; // @[Mux.scala 46:16:@11852.4]
  assign _T_14233 = 6'h1a == _T_10211_49; // @[Mux.scala 46:19:@11853.4]
  assign _T_14234 = _T_14233 ? _T_9260_25 : _T_14232; // @[Mux.scala 46:16:@11854.4]
  assign _T_14235 = 6'h19 == _T_10211_49; // @[Mux.scala 46:19:@11855.4]
  assign _T_14236 = _T_14235 ? _T_9260_24 : _T_14234; // @[Mux.scala 46:16:@11856.4]
  assign _T_14237 = 6'h18 == _T_10211_49; // @[Mux.scala 46:19:@11857.4]
  assign _T_14238 = _T_14237 ? _T_9260_23 : _T_14236; // @[Mux.scala 46:16:@11858.4]
  assign _T_14239 = 6'h17 == _T_10211_49; // @[Mux.scala 46:19:@11859.4]
  assign _T_14240 = _T_14239 ? _T_9260_22 : _T_14238; // @[Mux.scala 46:16:@11860.4]
  assign _T_14241 = 6'h16 == _T_10211_49; // @[Mux.scala 46:19:@11861.4]
  assign _T_14242 = _T_14241 ? _T_9260_21 : _T_14240; // @[Mux.scala 46:16:@11862.4]
  assign _T_14243 = 6'h15 == _T_10211_49; // @[Mux.scala 46:19:@11863.4]
  assign _T_14244 = _T_14243 ? _T_9260_20 : _T_14242; // @[Mux.scala 46:16:@11864.4]
  assign _T_14245 = 6'h14 == _T_10211_49; // @[Mux.scala 46:19:@11865.4]
  assign _T_14246 = _T_14245 ? _T_9260_19 : _T_14244; // @[Mux.scala 46:16:@11866.4]
  assign _T_14247 = 6'h13 == _T_10211_49; // @[Mux.scala 46:19:@11867.4]
  assign _T_14248 = _T_14247 ? _T_9260_18 : _T_14246; // @[Mux.scala 46:16:@11868.4]
  assign _T_14249 = 6'h12 == _T_10211_49; // @[Mux.scala 46:19:@11869.4]
  assign _T_14250 = _T_14249 ? _T_9260_17 : _T_14248; // @[Mux.scala 46:16:@11870.4]
  assign _T_14251 = 6'h11 == _T_10211_49; // @[Mux.scala 46:19:@11871.4]
  assign _T_14252 = _T_14251 ? _T_9260_16 : _T_14250; // @[Mux.scala 46:16:@11872.4]
  assign _T_14253 = 6'h10 == _T_10211_49; // @[Mux.scala 46:19:@11873.4]
  assign _T_14254 = _T_14253 ? _T_9260_15 : _T_14252; // @[Mux.scala 46:16:@11874.4]
  assign _T_14255 = 6'hf == _T_10211_49; // @[Mux.scala 46:19:@11875.4]
  assign _T_14256 = _T_14255 ? _T_9260_14 : _T_14254; // @[Mux.scala 46:16:@11876.4]
  assign _T_14257 = 6'he == _T_10211_49; // @[Mux.scala 46:19:@11877.4]
  assign _T_14258 = _T_14257 ? _T_9260_13 : _T_14256; // @[Mux.scala 46:16:@11878.4]
  assign _T_14259 = 6'hd == _T_10211_49; // @[Mux.scala 46:19:@11879.4]
  assign _T_14260 = _T_14259 ? _T_9260_12 : _T_14258; // @[Mux.scala 46:16:@11880.4]
  assign _T_14261 = 6'hc == _T_10211_49; // @[Mux.scala 46:19:@11881.4]
  assign _T_14262 = _T_14261 ? _T_9260_11 : _T_14260; // @[Mux.scala 46:16:@11882.4]
  assign _T_14263 = 6'hb == _T_10211_49; // @[Mux.scala 46:19:@11883.4]
  assign _T_14264 = _T_14263 ? _T_9260_10 : _T_14262; // @[Mux.scala 46:16:@11884.4]
  assign _T_14265 = 6'ha == _T_10211_49; // @[Mux.scala 46:19:@11885.4]
  assign _T_14266 = _T_14265 ? _T_9260_9 : _T_14264; // @[Mux.scala 46:16:@11886.4]
  assign _T_14267 = 6'h9 == _T_10211_49; // @[Mux.scala 46:19:@11887.4]
  assign _T_14268 = _T_14267 ? _T_9260_8 : _T_14266; // @[Mux.scala 46:16:@11888.4]
  assign _T_14269 = 6'h8 == _T_10211_49; // @[Mux.scala 46:19:@11889.4]
  assign _T_14270 = _T_14269 ? _T_9260_7 : _T_14268; // @[Mux.scala 46:16:@11890.4]
  assign _T_14271 = 6'h7 == _T_10211_49; // @[Mux.scala 46:19:@11891.4]
  assign _T_14272 = _T_14271 ? _T_9260_6 : _T_14270; // @[Mux.scala 46:16:@11892.4]
  assign _T_14273 = 6'h6 == _T_10211_49; // @[Mux.scala 46:19:@11893.4]
  assign _T_14274 = _T_14273 ? _T_9260_5 : _T_14272; // @[Mux.scala 46:16:@11894.4]
  assign _T_14275 = 6'h5 == _T_10211_49; // @[Mux.scala 46:19:@11895.4]
  assign _T_14276 = _T_14275 ? _T_9260_4 : _T_14274; // @[Mux.scala 46:16:@11896.4]
  assign _T_14277 = 6'h4 == _T_10211_49; // @[Mux.scala 46:19:@11897.4]
  assign _T_14278 = _T_14277 ? _T_9260_3 : _T_14276; // @[Mux.scala 46:16:@11898.4]
  assign _T_14279 = 6'h3 == _T_10211_49; // @[Mux.scala 46:19:@11899.4]
  assign _T_14280 = _T_14279 ? _T_9260_2 : _T_14278; // @[Mux.scala 46:16:@11900.4]
  assign _T_14281 = 6'h2 == _T_10211_49; // @[Mux.scala 46:19:@11901.4]
  assign _T_14282 = _T_14281 ? _T_9260_1 : _T_14280; // @[Mux.scala 46:16:@11902.4]
  assign _T_14283 = 6'h1 == _T_10211_49; // @[Mux.scala 46:19:@11903.4]
  assign _T_14284 = _T_14283 ? _T_9260_0 : _T_14282; // @[Mux.scala 46:16:@11904.4]
  assign _T_14337 = 6'h33 == _T_10211_50; // @[Mux.scala 46:19:@11906.4]
  assign _T_14338 = _T_14337 ? _T_9260_50 : 8'h0; // @[Mux.scala 46:16:@11907.4]
  assign _T_14339 = 6'h32 == _T_10211_50; // @[Mux.scala 46:19:@11908.4]
  assign _T_14340 = _T_14339 ? _T_9260_49 : _T_14338; // @[Mux.scala 46:16:@11909.4]
  assign _T_14341 = 6'h31 == _T_10211_50; // @[Mux.scala 46:19:@11910.4]
  assign _T_14342 = _T_14341 ? _T_9260_48 : _T_14340; // @[Mux.scala 46:16:@11911.4]
  assign _T_14343 = 6'h30 == _T_10211_50; // @[Mux.scala 46:19:@11912.4]
  assign _T_14344 = _T_14343 ? _T_9260_47 : _T_14342; // @[Mux.scala 46:16:@11913.4]
  assign _T_14345 = 6'h2f == _T_10211_50; // @[Mux.scala 46:19:@11914.4]
  assign _T_14346 = _T_14345 ? _T_9260_46 : _T_14344; // @[Mux.scala 46:16:@11915.4]
  assign _T_14347 = 6'h2e == _T_10211_50; // @[Mux.scala 46:19:@11916.4]
  assign _T_14348 = _T_14347 ? _T_9260_45 : _T_14346; // @[Mux.scala 46:16:@11917.4]
  assign _T_14349 = 6'h2d == _T_10211_50; // @[Mux.scala 46:19:@11918.4]
  assign _T_14350 = _T_14349 ? _T_9260_44 : _T_14348; // @[Mux.scala 46:16:@11919.4]
  assign _T_14351 = 6'h2c == _T_10211_50; // @[Mux.scala 46:19:@11920.4]
  assign _T_14352 = _T_14351 ? _T_9260_43 : _T_14350; // @[Mux.scala 46:16:@11921.4]
  assign _T_14353 = 6'h2b == _T_10211_50; // @[Mux.scala 46:19:@11922.4]
  assign _T_14354 = _T_14353 ? _T_9260_42 : _T_14352; // @[Mux.scala 46:16:@11923.4]
  assign _T_14355 = 6'h2a == _T_10211_50; // @[Mux.scala 46:19:@11924.4]
  assign _T_14356 = _T_14355 ? _T_9260_41 : _T_14354; // @[Mux.scala 46:16:@11925.4]
  assign _T_14357 = 6'h29 == _T_10211_50; // @[Mux.scala 46:19:@11926.4]
  assign _T_14358 = _T_14357 ? _T_9260_40 : _T_14356; // @[Mux.scala 46:16:@11927.4]
  assign _T_14359 = 6'h28 == _T_10211_50; // @[Mux.scala 46:19:@11928.4]
  assign _T_14360 = _T_14359 ? _T_9260_39 : _T_14358; // @[Mux.scala 46:16:@11929.4]
  assign _T_14361 = 6'h27 == _T_10211_50; // @[Mux.scala 46:19:@11930.4]
  assign _T_14362 = _T_14361 ? _T_9260_38 : _T_14360; // @[Mux.scala 46:16:@11931.4]
  assign _T_14363 = 6'h26 == _T_10211_50; // @[Mux.scala 46:19:@11932.4]
  assign _T_14364 = _T_14363 ? _T_9260_37 : _T_14362; // @[Mux.scala 46:16:@11933.4]
  assign _T_14365 = 6'h25 == _T_10211_50; // @[Mux.scala 46:19:@11934.4]
  assign _T_14366 = _T_14365 ? _T_9260_36 : _T_14364; // @[Mux.scala 46:16:@11935.4]
  assign _T_14367 = 6'h24 == _T_10211_50; // @[Mux.scala 46:19:@11936.4]
  assign _T_14368 = _T_14367 ? _T_9260_35 : _T_14366; // @[Mux.scala 46:16:@11937.4]
  assign _T_14369 = 6'h23 == _T_10211_50; // @[Mux.scala 46:19:@11938.4]
  assign _T_14370 = _T_14369 ? _T_9260_34 : _T_14368; // @[Mux.scala 46:16:@11939.4]
  assign _T_14371 = 6'h22 == _T_10211_50; // @[Mux.scala 46:19:@11940.4]
  assign _T_14372 = _T_14371 ? _T_9260_33 : _T_14370; // @[Mux.scala 46:16:@11941.4]
  assign _T_14373 = 6'h21 == _T_10211_50; // @[Mux.scala 46:19:@11942.4]
  assign _T_14374 = _T_14373 ? _T_9260_32 : _T_14372; // @[Mux.scala 46:16:@11943.4]
  assign _T_14375 = 6'h20 == _T_10211_50; // @[Mux.scala 46:19:@11944.4]
  assign _T_14376 = _T_14375 ? _T_9260_31 : _T_14374; // @[Mux.scala 46:16:@11945.4]
  assign _T_14377 = 6'h1f == _T_10211_50; // @[Mux.scala 46:19:@11946.4]
  assign _T_14378 = _T_14377 ? _T_9260_30 : _T_14376; // @[Mux.scala 46:16:@11947.4]
  assign _T_14379 = 6'h1e == _T_10211_50; // @[Mux.scala 46:19:@11948.4]
  assign _T_14380 = _T_14379 ? _T_9260_29 : _T_14378; // @[Mux.scala 46:16:@11949.4]
  assign _T_14381 = 6'h1d == _T_10211_50; // @[Mux.scala 46:19:@11950.4]
  assign _T_14382 = _T_14381 ? _T_9260_28 : _T_14380; // @[Mux.scala 46:16:@11951.4]
  assign _T_14383 = 6'h1c == _T_10211_50; // @[Mux.scala 46:19:@11952.4]
  assign _T_14384 = _T_14383 ? _T_9260_27 : _T_14382; // @[Mux.scala 46:16:@11953.4]
  assign _T_14385 = 6'h1b == _T_10211_50; // @[Mux.scala 46:19:@11954.4]
  assign _T_14386 = _T_14385 ? _T_9260_26 : _T_14384; // @[Mux.scala 46:16:@11955.4]
  assign _T_14387 = 6'h1a == _T_10211_50; // @[Mux.scala 46:19:@11956.4]
  assign _T_14388 = _T_14387 ? _T_9260_25 : _T_14386; // @[Mux.scala 46:16:@11957.4]
  assign _T_14389 = 6'h19 == _T_10211_50; // @[Mux.scala 46:19:@11958.4]
  assign _T_14390 = _T_14389 ? _T_9260_24 : _T_14388; // @[Mux.scala 46:16:@11959.4]
  assign _T_14391 = 6'h18 == _T_10211_50; // @[Mux.scala 46:19:@11960.4]
  assign _T_14392 = _T_14391 ? _T_9260_23 : _T_14390; // @[Mux.scala 46:16:@11961.4]
  assign _T_14393 = 6'h17 == _T_10211_50; // @[Mux.scala 46:19:@11962.4]
  assign _T_14394 = _T_14393 ? _T_9260_22 : _T_14392; // @[Mux.scala 46:16:@11963.4]
  assign _T_14395 = 6'h16 == _T_10211_50; // @[Mux.scala 46:19:@11964.4]
  assign _T_14396 = _T_14395 ? _T_9260_21 : _T_14394; // @[Mux.scala 46:16:@11965.4]
  assign _T_14397 = 6'h15 == _T_10211_50; // @[Mux.scala 46:19:@11966.4]
  assign _T_14398 = _T_14397 ? _T_9260_20 : _T_14396; // @[Mux.scala 46:16:@11967.4]
  assign _T_14399 = 6'h14 == _T_10211_50; // @[Mux.scala 46:19:@11968.4]
  assign _T_14400 = _T_14399 ? _T_9260_19 : _T_14398; // @[Mux.scala 46:16:@11969.4]
  assign _T_14401 = 6'h13 == _T_10211_50; // @[Mux.scala 46:19:@11970.4]
  assign _T_14402 = _T_14401 ? _T_9260_18 : _T_14400; // @[Mux.scala 46:16:@11971.4]
  assign _T_14403 = 6'h12 == _T_10211_50; // @[Mux.scala 46:19:@11972.4]
  assign _T_14404 = _T_14403 ? _T_9260_17 : _T_14402; // @[Mux.scala 46:16:@11973.4]
  assign _T_14405 = 6'h11 == _T_10211_50; // @[Mux.scala 46:19:@11974.4]
  assign _T_14406 = _T_14405 ? _T_9260_16 : _T_14404; // @[Mux.scala 46:16:@11975.4]
  assign _T_14407 = 6'h10 == _T_10211_50; // @[Mux.scala 46:19:@11976.4]
  assign _T_14408 = _T_14407 ? _T_9260_15 : _T_14406; // @[Mux.scala 46:16:@11977.4]
  assign _T_14409 = 6'hf == _T_10211_50; // @[Mux.scala 46:19:@11978.4]
  assign _T_14410 = _T_14409 ? _T_9260_14 : _T_14408; // @[Mux.scala 46:16:@11979.4]
  assign _T_14411 = 6'he == _T_10211_50; // @[Mux.scala 46:19:@11980.4]
  assign _T_14412 = _T_14411 ? _T_9260_13 : _T_14410; // @[Mux.scala 46:16:@11981.4]
  assign _T_14413 = 6'hd == _T_10211_50; // @[Mux.scala 46:19:@11982.4]
  assign _T_14414 = _T_14413 ? _T_9260_12 : _T_14412; // @[Mux.scala 46:16:@11983.4]
  assign _T_14415 = 6'hc == _T_10211_50; // @[Mux.scala 46:19:@11984.4]
  assign _T_14416 = _T_14415 ? _T_9260_11 : _T_14414; // @[Mux.scala 46:16:@11985.4]
  assign _T_14417 = 6'hb == _T_10211_50; // @[Mux.scala 46:19:@11986.4]
  assign _T_14418 = _T_14417 ? _T_9260_10 : _T_14416; // @[Mux.scala 46:16:@11987.4]
  assign _T_14419 = 6'ha == _T_10211_50; // @[Mux.scala 46:19:@11988.4]
  assign _T_14420 = _T_14419 ? _T_9260_9 : _T_14418; // @[Mux.scala 46:16:@11989.4]
  assign _T_14421 = 6'h9 == _T_10211_50; // @[Mux.scala 46:19:@11990.4]
  assign _T_14422 = _T_14421 ? _T_9260_8 : _T_14420; // @[Mux.scala 46:16:@11991.4]
  assign _T_14423 = 6'h8 == _T_10211_50; // @[Mux.scala 46:19:@11992.4]
  assign _T_14424 = _T_14423 ? _T_9260_7 : _T_14422; // @[Mux.scala 46:16:@11993.4]
  assign _T_14425 = 6'h7 == _T_10211_50; // @[Mux.scala 46:19:@11994.4]
  assign _T_14426 = _T_14425 ? _T_9260_6 : _T_14424; // @[Mux.scala 46:16:@11995.4]
  assign _T_14427 = 6'h6 == _T_10211_50; // @[Mux.scala 46:19:@11996.4]
  assign _T_14428 = _T_14427 ? _T_9260_5 : _T_14426; // @[Mux.scala 46:16:@11997.4]
  assign _T_14429 = 6'h5 == _T_10211_50; // @[Mux.scala 46:19:@11998.4]
  assign _T_14430 = _T_14429 ? _T_9260_4 : _T_14428; // @[Mux.scala 46:16:@11999.4]
  assign _T_14431 = 6'h4 == _T_10211_50; // @[Mux.scala 46:19:@12000.4]
  assign _T_14432 = _T_14431 ? _T_9260_3 : _T_14430; // @[Mux.scala 46:16:@12001.4]
  assign _T_14433 = 6'h3 == _T_10211_50; // @[Mux.scala 46:19:@12002.4]
  assign _T_14434 = _T_14433 ? _T_9260_2 : _T_14432; // @[Mux.scala 46:16:@12003.4]
  assign _T_14435 = 6'h2 == _T_10211_50; // @[Mux.scala 46:19:@12004.4]
  assign _T_14436 = _T_14435 ? _T_9260_1 : _T_14434; // @[Mux.scala 46:16:@12005.4]
  assign _T_14437 = 6'h1 == _T_10211_50; // @[Mux.scala 46:19:@12006.4]
  assign _T_14438 = _T_14437 ? _T_9260_0 : _T_14436; // @[Mux.scala 46:16:@12007.4]
  assign _T_14492 = 6'h34 == _T_10211_51; // @[Mux.scala 46:19:@12009.4]
  assign _T_14493 = _T_14492 ? _T_9260_51 : 8'h0; // @[Mux.scala 46:16:@12010.4]
  assign _T_14494 = 6'h33 == _T_10211_51; // @[Mux.scala 46:19:@12011.4]
  assign _T_14495 = _T_14494 ? _T_9260_50 : _T_14493; // @[Mux.scala 46:16:@12012.4]
  assign _T_14496 = 6'h32 == _T_10211_51; // @[Mux.scala 46:19:@12013.4]
  assign _T_14497 = _T_14496 ? _T_9260_49 : _T_14495; // @[Mux.scala 46:16:@12014.4]
  assign _T_14498 = 6'h31 == _T_10211_51; // @[Mux.scala 46:19:@12015.4]
  assign _T_14499 = _T_14498 ? _T_9260_48 : _T_14497; // @[Mux.scala 46:16:@12016.4]
  assign _T_14500 = 6'h30 == _T_10211_51; // @[Mux.scala 46:19:@12017.4]
  assign _T_14501 = _T_14500 ? _T_9260_47 : _T_14499; // @[Mux.scala 46:16:@12018.4]
  assign _T_14502 = 6'h2f == _T_10211_51; // @[Mux.scala 46:19:@12019.4]
  assign _T_14503 = _T_14502 ? _T_9260_46 : _T_14501; // @[Mux.scala 46:16:@12020.4]
  assign _T_14504 = 6'h2e == _T_10211_51; // @[Mux.scala 46:19:@12021.4]
  assign _T_14505 = _T_14504 ? _T_9260_45 : _T_14503; // @[Mux.scala 46:16:@12022.4]
  assign _T_14506 = 6'h2d == _T_10211_51; // @[Mux.scala 46:19:@12023.4]
  assign _T_14507 = _T_14506 ? _T_9260_44 : _T_14505; // @[Mux.scala 46:16:@12024.4]
  assign _T_14508 = 6'h2c == _T_10211_51; // @[Mux.scala 46:19:@12025.4]
  assign _T_14509 = _T_14508 ? _T_9260_43 : _T_14507; // @[Mux.scala 46:16:@12026.4]
  assign _T_14510 = 6'h2b == _T_10211_51; // @[Mux.scala 46:19:@12027.4]
  assign _T_14511 = _T_14510 ? _T_9260_42 : _T_14509; // @[Mux.scala 46:16:@12028.4]
  assign _T_14512 = 6'h2a == _T_10211_51; // @[Mux.scala 46:19:@12029.4]
  assign _T_14513 = _T_14512 ? _T_9260_41 : _T_14511; // @[Mux.scala 46:16:@12030.4]
  assign _T_14514 = 6'h29 == _T_10211_51; // @[Mux.scala 46:19:@12031.4]
  assign _T_14515 = _T_14514 ? _T_9260_40 : _T_14513; // @[Mux.scala 46:16:@12032.4]
  assign _T_14516 = 6'h28 == _T_10211_51; // @[Mux.scala 46:19:@12033.4]
  assign _T_14517 = _T_14516 ? _T_9260_39 : _T_14515; // @[Mux.scala 46:16:@12034.4]
  assign _T_14518 = 6'h27 == _T_10211_51; // @[Mux.scala 46:19:@12035.4]
  assign _T_14519 = _T_14518 ? _T_9260_38 : _T_14517; // @[Mux.scala 46:16:@12036.4]
  assign _T_14520 = 6'h26 == _T_10211_51; // @[Mux.scala 46:19:@12037.4]
  assign _T_14521 = _T_14520 ? _T_9260_37 : _T_14519; // @[Mux.scala 46:16:@12038.4]
  assign _T_14522 = 6'h25 == _T_10211_51; // @[Mux.scala 46:19:@12039.4]
  assign _T_14523 = _T_14522 ? _T_9260_36 : _T_14521; // @[Mux.scala 46:16:@12040.4]
  assign _T_14524 = 6'h24 == _T_10211_51; // @[Mux.scala 46:19:@12041.4]
  assign _T_14525 = _T_14524 ? _T_9260_35 : _T_14523; // @[Mux.scala 46:16:@12042.4]
  assign _T_14526 = 6'h23 == _T_10211_51; // @[Mux.scala 46:19:@12043.4]
  assign _T_14527 = _T_14526 ? _T_9260_34 : _T_14525; // @[Mux.scala 46:16:@12044.4]
  assign _T_14528 = 6'h22 == _T_10211_51; // @[Mux.scala 46:19:@12045.4]
  assign _T_14529 = _T_14528 ? _T_9260_33 : _T_14527; // @[Mux.scala 46:16:@12046.4]
  assign _T_14530 = 6'h21 == _T_10211_51; // @[Mux.scala 46:19:@12047.4]
  assign _T_14531 = _T_14530 ? _T_9260_32 : _T_14529; // @[Mux.scala 46:16:@12048.4]
  assign _T_14532 = 6'h20 == _T_10211_51; // @[Mux.scala 46:19:@12049.4]
  assign _T_14533 = _T_14532 ? _T_9260_31 : _T_14531; // @[Mux.scala 46:16:@12050.4]
  assign _T_14534 = 6'h1f == _T_10211_51; // @[Mux.scala 46:19:@12051.4]
  assign _T_14535 = _T_14534 ? _T_9260_30 : _T_14533; // @[Mux.scala 46:16:@12052.4]
  assign _T_14536 = 6'h1e == _T_10211_51; // @[Mux.scala 46:19:@12053.4]
  assign _T_14537 = _T_14536 ? _T_9260_29 : _T_14535; // @[Mux.scala 46:16:@12054.4]
  assign _T_14538 = 6'h1d == _T_10211_51; // @[Mux.scala 46:19:@12055.4]
  assign _T_14539 = _T_14538 ? _T_9260_28 : _T_14537; // @[Mux.scala 46:16:@12056.4]
  assign _T_14540 = 6'h1c == _T_10211_51; // @[Mux.scala 46:19:@12057.4]
  assign _T_14541 = _T_14540 ? _T_9260_27 : _T_14539; // @[Mux.scala 46:16:@12058.4]
  assign _T_14542 = 6'h1b == _T_10211_51; // @[Mux.scala 46:19:@12059.4]
  assign _T_14543 = _T_14542 ? _T_9260_26 : _T_14541; // @[Mux.scala 46:16:@12060.4]
  assign _T_14544 = 6'h1a == _T_10211_51; // @[Mux.scala 46:19:@12061.4]
  assign _T_14545 = _T_14544 ? _T_9260_25 : _T_14543; // @[Mux.scala 46:16:@12062.4]
  assign _T_14546 = 6'h19 == _T_10211_51; // @[Mux.scala 46:19:@12063.4]
  assign _T_14547 = _T_14546 ? _T_9260_24 : _T_14545; // @[Mux.scala 46:16:@12064.4]
  assign _T_14548 = 6'h18 == _T_10211_51; // @[Mux.scala 46:19:@12065.4]
  assign _T_14549 = _T_14548 ? _T_9260_23 : _T_14547; // @[Mux.scala 46:16:@12066.4]
  assign _T_14550 = 6'h17 == _T_10211_51; // @[Mux.scala 46:19:@12067.4]
  assign _T_14551 = _T_14550 ? _T_9260_22 : _T_14549; // @[Mux.scala 46:16:@12068.4]
  assign _T_14552 = 6'h16 == _T_10211_51; // @[Mux.scala 46:19:@12069.4]
  assign _T_14553 = _T_14552 ? _T_9260_21 : _T_14551; // @[Mux.scala 46:16:@12070.4]
  assign _T_14554 = 6'h15 == _T_10211_51; // @[Mux.scala 46:19:@12071.4]
  assign _T_14555 = _T_14554 ? _T_9260_20 : _T_14553; // @[Mux.scala 46:16:@12072.4]
  assign _T_14556 = 6'h14 == _T_10211_51; // @[Mux.scala 46:19:@12073.4]
  assign _T_14557 = _T_14556 ? _T_9260_19 : _T_14555; // @[Mux.scala 46:16:@12074.4]
  assign _T_14558 = 6'h13 == _T_10211_51; // @[Mux.scala 46:19:@12075.4]
  assign _T_14559 = _T_14558 ? _T_9260_18 : _T_14557; // @[Mux.scala 46:16:@12076.4]
  assign _T_14560 = 6'h12 == _T_10211_51; // @[Mux.scala 46:19:@12077.4]
  assign _T_14561 = _T_14560 ? _T_9260_17 : _T_14559; // @[Mux.scala 46:16:@12078.4]
  assign _T_14562 = 6'h11 == _T_10211_51; // @[Mux.scala 46:19:@12079.4]
  assign _T_14563 = _T_14562 ? _T_9260_16 : _T_14561; // @[Mux.scala 46:16:@12080.4]
  assign _T_14564 = 6'h10 == _T_10211_51; // @[Mux.scala 46:19:@12081.4]
  assign _T_14565 = _T_14564 ? _T_9260_15 : _T_14563; // @[Mux.scala 46:16:@12082.4]
  assign _T_14566 = 6'hf == _T_10211_51; // @[Mux.scala 46:19:@12083.4]
  assign _T_14567 = _T_14566 ? _T_9260_14 : _T_14565; // @[Mux.scala 46:16:@12084.4]
  assign _T_14568 = 6'he == _T_10211_51; // @[Mux.scala 46:19:@12085.4]
  assign _T_14569 = _T_14568 ? _T_9260_13 : _T_14567; // @[Mux.scala 46:16:@12086.4]
  assign _T_14570 = 6'hd == _T_10211_51; // @[Mux.scala 46:19:@12087.4]
  assign _T_14571 = _T_14570 ? _T_9260_12 : _T_14569; // @[Mux.scala 46:16:@12088.4]
  assign _T_14572 = 6'hc == _T_10211_51; // @[Mux.scala 46:19:@12089.4]
  assign _T_14573 = _T_14572 ? _T_9260_11 : _T_14571; // @[Mux.scala 46:16:@12090.4]
  assign _T_14574 = 6'hb == _T_10211_51; // @[Mux.scala 46:19:@12091.4]
  assign _T_14575 = _T_14574 ? _T_9260_10 : _T_14573; // @[Mux.scala 46:16:@12092.4]
  assign _T_14576 = 6'ha == _T_10211_51; // @[Mux.scala 46:19:@12093.4]
  assign _T_14577 = _T_14576 ? _T_9260_9 : _T_14575; // @[Mux.scala 46:16:@12094.4]
  assign _T_14578 = 6'h9 == _T_10211_51; // @[Mux.scala 46:19:@12095.4]
  assign _T_14579 = _T_14578 ? _T_9260_8 : _T_14577; // @[Mux.scala 46:16:@12096.4]
  assign _T_14580 = 6'h8 == _T_10211_51; // @[Mux.scala 46:19:@12097.4]
  assign _T_14581 = _T_14580 ? _T_9260_7 : _T_14579; // @[Mux.scala 46:16:@12098.4]
  assign _T_14582 = 6'h7 == _T_10211_51; // @[Mux.scala 46:19:@12099.4]
  assign _T_14583 = _T_14582 ? _T_9260_6 : _T_14581; // @[Mux.scala 46:16:@12100.4]
  assign _T_14584 = 6'h6 == _T_10211_51; // @[Mux.scala 46:19:@12101.4]
  assign _T_14585 = _T_14584 ? _T_9260_5 : _T_14583; // @[Mux.scala 46:16:@12102.4]
  assign _T_14586 = 6'h5 == _T_10211_51; // @[Mux.scala 46:19:@12103.4]
  assign _T_14587 = _T_14586 ? _T_9260_4 : _T_14585; // @[Mux.scala 46:16:@12104.4]
  assign _T_14588 = 6'h4 == _T_10211_51; // @[Mux.scala 46:19:@12105.4]
  assign _T_14589 = _T_14588 ? _T_9260_3 : _T_14587; // @[Mux.scala 46:16:@12106.4]
  assign _T_14590 = 6'h3 == _T_10211_51; // @[Mux.scala 46:19:@12107.4]
  assign _T_14591 = _T_14590 ? _T_9260_2 : _T_14589; // @[Mux.scala 46:16:@12108.4]
  assign _T_14592 = 6'h2 == _T_10211_51; // @[Mux.scala 46:19:@12109.4]
  assign _T_14593 = _T_14592 ? _T_9260_1 : _T_14591; // @[Mux.scala 46:16:@12110.4]
  assign _T_14594 = 6'h1 == _T_10211_51; // @[Mux.scala 46:19:@12111.4]
  assign _T_14595 = _T_14594 ? _T_9260_0 : _T_14593; // @[Mux.scala 46:16:@12112.4]
  assign _T_14650 = 6'h35 == _T_10211_52; // @[Mux.scala 46:19:@12114.4]
  assign _T_14651 = _T_14650 ? _T_9260_52 : 8'h0; // @[Mux.scala 46:16:@12115.4]
  assign _T_14652 = 6'h34 == _T_10211_52; // @[Mux.scala 46:19:@12116.4]
  assign _T_14653 = _T_14652 ? _T_9260_51 : _T_14651; // @[Mux.scala 46:16:@12117.4]
  assign _T_14654 = 6'h33 == _T_10211_52; // @[Mux.scala 46:19:@12118.4]
  assign _T_14655 = _T_14654 ? _T_9260_50 : _T_14653; // @[Mux.scala 46:16:@12119.4]
  assign _T_14656 = 6'h32 == _T_10211_52; // @[Mux.scala 46:19:@12120.4]
  assign _T_14657 = _T_14656 ? _T_9260_49 : _T_14655; // @[Mux.scala 46:16:@12121.4]
  assign _T_14658 = 6'h31 == _T_10211_52; // @[Mux.scala 46:19:@12122.4]
  assign _T_14659 = _T_14658 ? _T_9260_48 : _T_14657; // @[Mux.scala 46:16:@12123.4]
  assign _T_14660 = 6'h30 == _T_10211_52; // @[Mux.scala 46:19:@12124.4]
  assign _T_14661 = _T_14660 ? _T_9260_47 : _T_14659; // @[Mux.scala 46:16:@12125.4]
  assign _T_14662 = 6'h2f == _T_10211_52; // @[Mux.scala 46:19:@12126.4]
  assign _T_14663 = _T_14662 ? _T_9260_46 : _T_14661; // @[Mux.scala 46:16:@12127.4]
  assign _T_14664 = 6'h2e == _T_10211_52; // @[Mux.scala 46:19:@12128.4]
  assign _T_14665 = _T_14664 ? _T_9260_45 : _T_14663; // @[Mux.scala 46:16:@12129.4]
  assign _T_14666 = 6'h2d == _T_10211_52; // @[Mux.scala 46:19:@12130.4]
  assign _T_14667 = _T_14666 ? _T_9260_44 : _T_14665; // @[Mux.scala 46:16:@12131.4]
  assign _T_14668 = 6'h2c == _T_10211_52; // @[Mux.scala 46:19:@12132.4]
  assign _T_14669 = _T_14668 ? _T_9260_43 : _T_14667; // @[Mux.scala 46:16:@12133.4]
  assign _T_14670 = 6'h2b == _T_10211_52; // @[Mux.scala 46:19:@12134.4]
  assign _T_14671 = _T_14670 ? _T_9260_42 : _T_14669; // @[Mux.scala 46:16:@12135.4]
  assign _T_14672 = 6'h2a == _T_10211_52; // @[Mux.scala 46:19:@12136.4]
  assign _T_14673 = _T_14672 ? _T_9260_41 : _T_14671; // @[Mux.scala 46:16:@12137.4]
  assign _T_14674 = 6'h29 == _T_10211_52; // @[Mux.scala 46:19:@12138.4]
  assign _T_14675 = _T_14674 ? _T_9260_40 : _T_14673; // @[Mux.scala 46:16:@12139.4]
  assign _T_14676 = 6'h28 == _T_10211_52; // @[Mux.scala 46:19:@12140.4]
  assign _T_14677 = _T_14676 ? _T_9260_39 : _T_14675; // @[Mux.scala 46:16:@12141.4]
  assign _T_14678 = 6'h27 == _T_10211_52; // @[Mux.scala 46:19:@12142.4]
  assign _T_14679 = _T_14678 ? _T_9260_38 : _T_14677; // @[Mux.scala 46:16:@12143.4]
  assign _T_14680 = 6'h26 == _T_10211_52; // @[Mux.scala 46:19:@12144.4]
  assign _T_14681 = _T_14680 ? _T_9260_37 : _T_14679; // @[Mux.scala 46:16:@12145.4]
  assign _T_14682 = 6'h25 == _T_10211_52; // @[Mux.scala 46:19:@12146.4]
  assign _T_14683 = _T_14682 ? _T_9260_36 : _T_14681; // @[Mux.scala 46:16:@12147.4]
  assign _T_14684 = 6'h24 == _T_10211_52; // @[Mux.scala 46:19:@12148.4]
  assign _T_14685 = _T_14684 ? _T_9260_35 : _T_14683; // @[Mux.scala 46:16:@12149.4]
  assign _T_14686 = 6'h23 == _T_10211_52; // @[Mux.scala 46:19:@12150.4]
  assign _T_14687 = _T_14686 ? _T_9260_34 : _T_14685; // @[Mux.scala 46:16:@12151.4]
  assign _T_14688 = 6'h22 == _T_10211_52; // @[Mux.scala 46:19:@12152.4]
  assign _T_14689 = _T_14688 ? _T_9260_33 : _T_14687; // @[Mux.scala 46:16:@12153.4]
  assign _T_14690 = 6'h21 == _T_10211_52; // @[Mux.scala 46:19:@12154.4]
  assign _T_14691 = _T_14690 ? _T_9260_32 : _T_14689; // @[Mux.scala 46:16:@12155.4]
  assign _T_14692 = 6'h20 == _T_10211_52; // @[Mux.scala 46:19:@12156.4]
  assign _T_14693 = _T_14692 ? _T_9260_31 : _T_14691; // @[Mux.scala 46:16:@12157.4]
  assign _T_14694 = 6'h1f == _T_10211_52; // @[Mux.scala 46:19:@12158.4]
  assign _T_14695 = _T_14694 ? _T_9260_30 : _T_14693; // @[Mux.scala 46:16:@12159.4]
  assign _T_14696 = 6'h1e == _T_10211_52; // @[Mux.scala 46:19:@12160.4]
  assign _T_14697 = _T_14696 ? _T_9260_29 : _T_14695; // @[Mux.scala 46:16:@12161.4]
  assign _T_14698 = 6'h1d == _T_10211_52; // @[Mux.scala 46:19:@12162.4]
  assign _T_14699 = _T_14698 ? _T_9260_28 : _T_14697; // @[Mux.scala 46:16:@12163.4]
  assign _T_14700 = 6'h1c == _T_10211_52; // @[Mux.scala 46:19:@12164.4]
  assign _T_14701 = _T_14700 ? _T_9260_27 : _T_14699; // @[Mux.scala 46:16:@12165.4]
  assign _T_14702 = 6'h1b == _T_10211_52; // @[Mux.scala 46:19:@12166.4]
  assign _T_14703 = _T_14702 ? _T_9260_26 : _T_14701; // @[Mux.scala 46:16:@12167.4]
  assign _T_14704 = 6'h1a == _T_10211_52; // @[Mux.scala 46:19:@12168.4]
  assign _T_14705 = _T_14704 ? _T_9260_25 : _T_14703; // @[Mux.scala 46:16:@12169.4]
  assign _T_14706 = 6'h19 == _T_10211_52; // @[Mux.scala 46:19:@12170.4]
  assign _T_14707 = _T_14706 ? _T_9260_24 : _T_14705; // @[Mux.scala 46:16:@12171.4]
  assign _T_14708 = 6'h18 == _T_10211_52; // @[Mux.scala 46:19:@12172.4]
  assign _T_14709 = _T_14708 ? _T_9260_23 : _T_14707; // @[Mux.scala 46:16:@12173.4]
  assign _T_14710 = 6'h17 == _T_10211_52; // @[Mux.scala 46:19:@12174.4]
  assign _T_14711 = _T_14710 ? _T_9260_22 : _T_14709; // @[Mux.scala 46:16:@12175.4]
  assign _T_14712 = 6'h16 == _T_10211_52; // @[Mux.scala 46:19:@12176.4]
  assign _T_14713 = _T_14712 ? _T_9260_21 : _T_14711; // @[Mux.scala 46:16:@12177.4]
  assign _T_14714 = 6'h15 == _T_10211_52; // @[Mux.scala 46:19:@12178.4]
  assign _T_14715 = _T_14714 ? _T_9260_20 : _T_14713; // @[Mux.scala 46:16:@12179.4]
  assign _T_14716 = 6'h14 == _T_10211_52; // @[Mux.scala 46:19:@12180.4]
  assign _T_14717 = _T_14716 ? _T_9260_19 : _T_14715; // @[Mux.scala 46:16:@12181.4]
  assign _T_14718 = 6'h13 == _T_10211_52; // @[Mux.scala 46:19:@12182.4]
  assign _T_14719 = _T_14718 ? _T_9260_18 : _T_14717; // @[Mux.scala 46:16:@12183.4]
  assign _T_14720 = 6'h12 == _T_10211_52; // @[Mux.scala 46:19:@12184.4]
  assign _T_14721 = _T_14720 ? _T_9260_17 : _T_14719; // @[Mux.scala 46:16:@12185.4]
  assign _T_14722 = 6'h11 == _T_10211_52; // @[Mux.scala 46:19:@12186.4]
  assign _T_14723 = _T_14722 ? _T_9260_16 : _T_14721; // @[Mux.scala 46:16:@12187.4]
  assign _T_14724 = 6'h10 == _T_10211_52; // @[Mux.scala 46:19:@12188.4]
  assign _T_14725 = _T_14724 ? _T_9260_15 : _T_14723; // @[Mux.scala 46:16:@12189.4]
  assign _T_14726 = 6'hf == _T_10211_52; // @[Mux.scala 46:19:@12190.4]
  assign _T_14727 = _T_14726 ? _T_9260_14 : _T_14725; // @[Mux.scala 46:16:@12191.4]
  assign _T_14728 = 6'he == _T_10211_52; // @[Mux.scala 46:19:@12192.4]
  assign _T_14729 = _T_14728 ? _T_9260_13 : _T_14727; // @[Mux.scala 46:16:@12193.4]
  assign _T_14730 = 6'hd == _T_10211_52; // @[Mux.scala 46:19:@12194.4]
  assign _T_14731 = _T_14730 ? _T_9260_12 : _T_14729; // @[Mux.scala 46:16:@12195.4]
  assign _T_14732 = 6'hc == _T_10211_52; // @[Mux.scala 46:19:@12196.4]
  assign _T_14733 = _T_14732 ? _T_9260_11 : _T_14731; // @[Mux.scala 46:16:@12197.4]
  assign _T_14734 = 6'hb == _T_10211_52; // @[Mux.scala 46:19:@12198.4]
  assign _T_14735 = _T_14734 ? _T_9260_10 : _T_14733; // @[Mux.scala 46:16:@12199.4]
  assign _T_14736 = 6'ha == _T_10211_52; // @[Mux.scala 46:19:@12200.4]
  assign _T_14737 = _T_14736 ? _T_9260_9 : _T_14735; // @[Mux.scala 46:16:@12201.4]
  assign _T_14738 = 6'h9 == _T_10211_52; // @[Mux.scala 46:19:@12202.4]
  assign _T_14739 = _T_14738 ? _T_9260_8 : _T_14737; // @[Mux.scala 46:16:@12203.4]
  assign _T_14740 = 6'h8 == _T_10211_52; // @[Mux.scala 46:19:@12204.4]
  assign _T_14741 = _T_14740 ? _T_9260_7 : _T_14739; // @[Mux.scala 46:16:@12205.4]
  assign _T_14742 = 6'h7 == _T_10211_52; // @[Mux.scala 46:19:@12206.4]
  assign _T_14743 = _T_14742 ? _T_9260_6 : _T_14741; // @[Mux.scala 46:16:@12207.4]
  assign _T_14744 = 6'h6 == _T_10211_52; // @[Mux.scala 46:19:@12208.4]
  assign _T_14745 = _T_14744 ? _T_9260_5 : _T_14743; // @[Mux.scala 46:16:@12209.4]
  assign _T_14746 = 6'h5 == _T_10211_52; // @[Mux.scala 46:19:@12210.4]
  assign _T_14747 = _T_14746 ? _T_9260_4 : _T_14745; // @[Mux.scala 46:16:@12211.4]
  assign _T_14748 = 6'h4 == _T_10211_52; // @[Mux.scala 46:19:@12212.4]
  assign _T_14749 = _T_14748 ? _T_9260_3 : _T_14747; // @[Mux.scala 46:16:@12213.4]
  assign _T_14750 = 6'h3 == _T_10211_52; // @[Mux.scala 46:19:@12214.4]
  assign _T_14751 = _T_14750 ? _T_9260_2 : _T_14749; // @[Mux.scala 46:16:@12215.4]
  assign _T_14752 = 6'h2 == _T_10211_52; // @[Mux.scala 46:19:@12216.4]
  assign _T_14753 = _T_14752 ? _T_9260_1 : _T_14751; // @[Mux.scala 46:16:@12217.4]
  assign _T_14754 = 6'h1 == _T_10211_52; // @[Mux.scala 46:19:@12218.4]
  assign _T_14755 = _T_14754 ? _T_9260_0 : _T_14753; // @[Mux.scala 46:16:@12219.4]
  assign _T_14811 = 6'h36 == _T_10211_53; // @[Mux.scala 46:19:@12221.4]
  assign _T_14812 = _T_14811 ? _T_9260_53 : 8'h0; // @[Mux.scala 46:16:@12222.4]
  assign _T_14813 = 6'h35 == _T_10211_53; // @[Mux.scala 46:19:@12223.4]
  assign _T_14814 = _T_14813 ? _T_9260_52 : _T_14812; // @[Mux.scala 46:16:@12224.4]
  assign _T_14815 = 6'h34 == _T_10211_53; // @[Mux.scala 46:19:@12225.4]
  assign _T_14816 = _T_14815 ? _T_9260_51 : _T_14814; // @[Mux.scala 46:16:@12226.4]
  assign _T_14817 = 6'h33 == _T_10211_53; // @[Mux.scala 46:19:@12227.4]
  assign _T_14818 = _T_14817 ? _T_9260_50 : _T_14816; // @[Mux.scala 46:16:@12228.4]
  assign _T_14819 = 6'h32 == _T_10211_53; // @[Mux.scala 46:19:@12229.4]
  assign _T_14820 = _T_14819 ? _T_9260_49 : _T_14818; // @[Mux.scala 46:16:@12230.4]
  assign _T_14821 = 6'h31 == _T_10211_53; // @[Mux.scala 46:19:@12231.4]
  assign _T_14822 = _T_14821 ? _T_9260_48 : _T_14820; // @[Mux.scala 46:16:@12232.4]
  assign _T_14823 = 6'h30 == _T_10211_53; // @[Mux.scala 46:19:@12233.4]
  assign _T_14824 = _T_14823 ? _T_9260_47 : _T_14822; // @[Mux.scala 46:16:@12234.4]
  assign _T_14825 = 6'h2f == _T_10211_53; // @[Mux.scala 46:19:@12235.4]
  assign _T_14826 = _T_14825 ? _T_9260_46 : _T_14824; // @[Mux.scala 46:16:@12236.4]
  assign _T_14827 = 6'h2e == _T_10211_53; // @[Mux.scala 46:19:@12237.4]
  assign _T_14828 = _T_14827 ? _T_9260_45 : _T_14826; // @[Mux.scala 46:16:@12238.4]
  assign _T_14829 = 6'h2d == _T_10211_53; // @[Mux.scala 46:19:@12239.4]
  assign _T_14830 = _T_14829 ? _T_9260_44 : _T_14828; // @[Mux.scala 46:16:@12240.4]
  assign _T_14831 = 6'h2c == _T_10211_53; // @[Mux.scala 46:19:@12241.4]
  assign _T_14832 = _T_14831 ? _T_9260_43 : _T_14830; // @[Mux.scala 46:16:@12242.4]
  assign _T_14833 = 6'h2b == _T_10211_53; // @[Mux.scala 46:19:@12243.4]
  assign _T_14834 = _T_14833 ? _T_9260_42 : _T_14832; // @[Mux.scala 46:16:@12244.4]
  assign _T_14835 = 6'h2a == _T_10211_53; // @[Mux.scala 46:19:@12245.4]
  assign _T_14836 = _T_14835 ? _T_9260_41 : _T_14834; // @[Mux.scala 46:16:@12246.4]
  assign _T_14837 = 6'h29 == _T_10211_53; // @[Mux.scala 46:19:@12247.4]
  assign _T_14838 = _T_14837 ? _T_9260_40 : _T_14836; // @[Mux.scala 46:16:@12248.4]
  assign _T_14839 = 6'h28 == _T_10211_53; // @[Mux.scala 46:19:@12249.4]
  assign _T_14840 = _T_14839 ? _T_9260_39 : _T_14838; // @[Mux.scala 46:16:@12250.4]
  assign _T_14841 = 6'h27 == _T_10211_53; // @[Mux.scala 46:19:@12251.4]
  assign _T_14842 = _T_14841 ? _T_9260_38 : _T_14840; // @[Mux.scala 46:16:@12252.4]
  assign _T_14843 = 6'h26 == _T_10211_53; // @[Mux.scala 46:19:@12253.4]
  assign _T_14844 = _T_14843 ? _T_9260_37 : _T_14842; // @[Mux.scala 46:16:@12254.4]
  assign _T_14845 = 6'h25 == _T_10211_53; // @[Mux.scala 46:19:@12255.4]
  assign _T_14846 = _T_14845 ? _T_9260_36 : _T_14844; // @[Mux.scala 46:16:@12256.4]
  assign _T_14847 = 6'h24 == _T_10211_53; // @[Mux.scala 46:19:@12257.4]
  assign _T_14848 = _T_14847 ? _T_9260_35 : _T_14846; // @[Mux.scala 46:16:@12258.4]
  assign _T_14849 = 6'h23 == _T_10211_53; // @[Mux.scala 46:19:@12259.4]
  assign _T_14850 = _T_14849 ? _T_9260_34 : _T_14848; // @[Mux.scala 46:16:@12260.4]
  assign _T_14851 = 6'h22 == _T_10211_53; // @[Mux.scala 46:19:@12261.4]
  assign _T_14852 = _T_14851 ? _T_9260_33 : _T_14850; // @[Mux.scala 46:16:@12262.4]
  assign _T_14853 = 6'h21 == _T_10211_53; // @[Mux.scala 46:19:@12263.4]
  assign _T_14854 = _T_14853 ? _T_9260_32 : _T_14852; // @[Mux.scala 46:16:@12264.4]
  assign _T_14855 = 6'h20 == _T_10211_53; // @[Mux.scala 46:19:@12265.4]
  assign _T_14856 = _T_14855 ? _T_9260_31 : _T_14854; // @[Mux.scala 46:16:@12266.4]
  assign _T_14857 = 6'h1f == _T_10211_53; // @[Mux.scala 46:19:@12267.4]
  assign _T_14858 = _T_14857 ? _T_9260_30 : _T_14856; // @[Mux.scala 46:16:@12268.4]
  assign _T_14859 = 6'h1e == _T_10211_53; // @[Mux.scala 46:19:@12269.4]
  assign _T_14860 = _T_14859 ? _T_9260_29 : _T_14858; // @[Mux.scala 46:16:@12270.4]
  assign _T_14861 = 6'h1d == _T_10211_53; // @[Mux.scala 46:19:@12271.4]
  assign _T_14862 = _T_14861 ? _T_9260_28 : _T_14860; // @[Mux.scala 46:16:@12272.4]
  assign _T_14863 = 6'h1c == _T_10211_53; // @[Mux.scala 46:19:@12273.4]
  assign _T_14864 = _T_14863 ? _T_9260_27 : _T_14862; // @[Mux.scala 46:16:@12274.4]
  assign _T_14865 = 6'h1b == _T_10211_53; // @[Mux.scala 46:19:@12275.4]
  assign _T_14866 = _T_14865 ? _T_9260_26 : _T_14864; // @[Mux.scala 46:16:@12276.4]
  assign _T_14867 = 6'h1a == _T_10211_53; // @[Mux.scala 46:19:@12277.4]
  assign _T_14868 = _T_14867 ? _T_9260_25 : _T_14866; // @[Mux.scala 46:16:@12278.4]
  assign _T_14869 = 6'h19 == _T_10211_53; // @[Mux.scala 46:19:@12279.4]
  assign _T_14870 = _T_14869 ? _T_9260_24 : _T_14868; // @[Mux.scala 46:16:@12280.4]
  assign _T_14871 = 6'h18 == _T_10211_53; // @[Mux.scala 46:19:@12281.4]
  assign _T_14872 = _T_14871 ? _T_9260_23 : _T_14870; // @[Mux.scala 46:16:@12282.4]
  assign _T_14873 = 6'h17 == _T_10211_53; // @[Mux.scala 46:19:@12283.4]
  assign _T_14874 = _T_14873 ? _T_9260_22 : _T_14872; // @[Mux.scala 46:16:@12284.4]
  assign _T_14875 = 6'h16 == _T_10211_53; // @[Mux.scala 46:19:@12285.4]
  assign _T_14876 = _T_14875 ? _T_9260_21 : _T_14874; // @[Mux.scala 46:16:@12286.4]
  assign _T_14877 = 6'h15 == _T_10211_53; // @[Mux.scala 46:19:@12287.4]
  assign _T_14878 = _T_14877 ? _T_9260_20 : _T_14876; // @[Mux.scala 46:16:@12288.4]
  assign _T_14879 = 6'h14 == _T_10211_53; // @[Mux.scala 46:19:@12289.4]
  assign _T_14880 = _T_14879 ? _T_9260_19 : _T_14878; // @[Mux.scala 46:16:@12290.4]
  assign _T_14881 = 6'h13 == _T_10211_53; // @[Mux.scala 46:19:@12291.4]
  assign _T_14882 = _T_14881 ? _T_9260_18 : _T_14880; // @[Mux.scala 46:16:@12292.4]
  assign _T_14883 = 6'h12 == _T_10211_53; // @[Mux.scala 46:19:@12293.4]
  assign _T_14884 = _T_14883 ? _T_9260_17 : _T_14882; // @[Mux.scala 46:16:@12294.4]
  assign _T_14885 = 6'h11 == _T_10211_53; // @[Mux.scala 46:19:@12295.4]
  assign _T_14886 = _T_14885 ? _T_9260_16 : _T_14884; // @[Mux.scala 46:16:@12296.4]
  assign _T_14887 = 6'h10 == _T_10211_53; // @[Mux.scala 46:19:@12297.4]
  assign _T_14888 = _T_14887 ? _T_9260_15 : _T_14886; // @[Mux.scala 46:16:@12298.4]
  assign _T_14889 = 6'hf == _T_10211_53; // @[Mux.scala 46:19:@12299.4]
  assign _T_14890 = _T_14889 ? _T_9260_14 : _T_14888; // @[Mux.scala 46:16:@12300.4]
  assign _T_14891 = 6'he == _T_10211_53; // @[Mux.scala 46:19:@12301.4]
  assign _T_14892 = _T_14891 ? _T_9260_13 : _T_14890; // @[Mux.scala 46:16:@12302.4]
  assign _T_14893 = 6'hd == _T_10211_53; // @[Mux.scala 46:19:@12303.4]
  assign _T_14894 = _T_14893 ? _T_9260_12 : _T_14892; // @[Mux.scala 46:16:@12304.4]
  assign _T_14895 = 6'hc == _T_10211_53; // @[Mux.scala 46:19:@12305.4]
  assign _T_14896 = _T_14895 ? _T_9260_11 : _T_14894; // @[Mux.scala 46:16:@12306.4]
  assign _T_14897 = 6'hb == _T_10211_53; // @[Mux.scala 46:19:@12307.4]
  assign _T_14898 = _T_14897 ? _T_9260_10 : _T_14896; // @[Mux.scala 46:16:@12308.4]
  assign _T_14899 = 6'ha == _T_10211_53; // @[Mux.scala 46:19:@12309.4]
  assign _T_14900 = _T_14899 ? _T_9260_9 : _T_14898; // @[Mux.scala 46:16:@12310.4]
  assign _T_14901 = 6'h9 == _T_10211_53; // @[Mux.scala 46:19:@12311.4]
  assign _T_14902 = _T_14901 ? _T_9260_8 : _T_14900; // @[Mux.scala 46:16:@12312.4]
  assign _T_14903 = 6'h8 == _T_10211_53; // @[Mux.scala 46:19:@12313.4]
  assign _T_14904 = _T_14903 ? _T_9260_7 : _T_14902; // @[Mux.scala 46:16:@12314.4]
  assign _T_14905 = 6'h7 == _T_10211_53; // @[Mux.scala 46:19:@12315.4]
  assign _T_14906 = _T_14905 ? _T_9260_6 : _T_14904; // @[Mux.scala 46:16:@12316.4]
  assign _T_14907 = 6'h6 == _T_10211_53; // @[Mux.scala 46:19:@12317.4]
  assign _T_14908 = _T_14907 ? _T_9260_5 : _T_14906; // @[Mux.scala 46:16:@12318.4]
  assign _T_14909 = 6'h5 == _T_10211_53; // @[Mux.scala 46:19:@12319.4]
  assign _T_14910 = _T_14909 ? _T_9260_4 : _T_14908; // @[Mux.scala 46:16:@12320.4]
  assign _T_14911 = 6'h4 == _T_10211_53; // @[Mux.scala 46:19:@12321.4]
  assign _T_14912 = _T_14911 ? _T_9260_3 : _T_14910; // @[Mux.scala 46:16:@12322.4]
  assign _T_14913 = 6'h3 == _T_10211_53; // @[Mux.scala 46:19:@12323.4]
  assign _T_14914 = _T_14913 ? _T_9260_2 : _T_14912; // @[Mux.scala 46:16:@12324.4]
  assign _T_14915 = 6'h2 == _T_10211_53; // @[Mux.scala 46:19:@12325.4]
  assign _T_14916 = _T_14915 ? _T_9260_1 : _T_14914; // @[Mux.scala 46:16:@12326.4]
  assign _T_14917 = 6'h1 == _T_10211_53; // @[Mux.scala 46:19:@12327.4]
  assign _T_14918 = _T_14917 ? _T_9260_0 : _T_14916; // @[Mux.scala 46:16:@12328.4]
  assign _T_14975 = 6'h37 == _T_10211_54; // @[Mux.scala 46:19:@12330.4]
  assign _T_14976 = _T_14975 ? _T_9260_54 : 8'h0; // @[Mux.scala 46:16:@12331.4]
  assign _T_14977 = 6'h36 == _T_10211_54; // @[Mux.scala 46:19:@12332.4]
  assign _T_14978 = _T_14977 ? _T_9260_53 : _T_14976; // @[Mux.scala 46:16:@12333.4]
  assign _T_14979 = 6'h35 == _T_10211_54; // @[Mux.scala 46:19:@12334.4]
  assign _T_14980 = _T_14979 ? _T_9260_52 : _T_14978; // @[Mux.scala 46:16:@12335.4]
  assign _T_14981 = 6'h34 == _T_10211_54; // @[Mux.scala 46:19:@12336.4]
  assign _T_14982 = _T_14981 ? _T_9260_51 : _T_14980; // @[Mux.scala 46:16:@12337.4]
  assign _T_14983 = 6'h33 == _T_10211_54; // @[Mux.scala 46:19:@12338.4]
  assign _T_14984 = _T_14983 ? _T_9260_50 : _T_14982; // @[Mux.scala 46:16:@12339.4]
  assign _T_14985 = 6'h32 == _T_10211_54; // @[Mux.scala 46:19:@12340.4]
  assign _T_14986 = _T_14985 ? _T_9260_49 : _T_14984; // @[Mux.scala 46:16:@12341.4]
  assign _T_14987 = 6'h31 == _T_10211_54; // @[Mux.scala 46:19:@12342.4]
  assign _T_14988 = _T_14987 ? _T_9260_48 : _T_14986; // @[Mux.scala 46:16:@12343.4]
  assign _T_14989 = 6'h30 == _T_10211_54; // @[Mux.scala 46:19:@12344.4]
  assign _T_14990 = _T_14989 ? _T_9260_47 : _T_14988; // @[Mux.scala 46:16:@12345.4]
  assign _T_14991 = 6'h2f == _T_10211_54; // @[Mux.scala 46:19:@12346.4]
  assign _T_14992 = _T_14991 ? _T_9260_46 : _T_14990; // @[Mux.scala 46:16:@12347.4]
  assign _T_14993 = 6'h2e == _T_10211_54; // @[Mux.scala 46:19:@12348.4]
  assign _T_14994 = _T_14993 ? _T_9260_45 : _T_14992; // @[Mux.scala 46:16:@12349.4]
  assign _T_14995 = 6'h2d == _T_10211_54; // @[Mux.scala 46:19:@12350.4]
  assign _T_14996 = _T_14995 ? _T_9260_44 : _T_14994; // @[Mux.scala 46:16:@12351.4]
  assign _T_14997 = 6'h2c == _T_10211_54; // @[Mux.scala 46:19:@12352.4]
  assign _T_14998 = _T_14997 ? _T_9260_43 : _T_14996; // @[Mux.scala 46:16:@12353.4]
  assign _T_14999 = 6'h2b == _T_10211_54; // @[Mux.scala 46:19:@12354.4]
  assign _T_15000 = _T_14999 ? _T_9260_42 : _T_14998; // @[Mux.scala 46:16:@12355.4]
  assign _T_15001 = 6'h2a == _T_10211_54; // @[Mux.scala 46:19:@12356.4]
  assign _T_15002 = _T_15001 ? _T_9260_41 : _T_15000; // @[Mux.scala 46:16:@12357.4]
  assign _T_15003 = 6'h29 == _T_10211_54; // @[Mux.scala 46:19:@12358.4]
  assign _T_15004 = _T_15003 ? _T_9260_40 : _T_15002; // @[Mux.scala 46:16:@12359.4]
  assign _T_15005 = 6'h28 == _T_10211_54; // @[Mux.scala 46:19:@12360.4]
  assign _T_15006 = _T_15005 ? _T_9260_39 : _T_15004; // @[Mux.scala 46:16:@12361.4]
  assign _T_15007 = 6'h27 == _T_10211_54; // @[Mux.scala 46:19:@12362.4]
  assign _T_15008 = _T_15007 ? _T_9260_38 : _T_15006; // @[Mux.scala 46:16:@12363.4]
  assign _T_15009 = 6'h26 == _T_10211_54; // @[Mux.scala 46:19:@12364.4]
  assign _T_15010 = _T_15009 ? _T_9260_37 : _T_15008; // @[Mux.scala 46:16:@12365.4]
  assign _T_15011 = 6'h25 == _T_10211_54; // @[Mux.scala 46:19:@12366.4]
  assign _T_15012 = _T_15011 ? _T_9260_36 : _T_15010; // @[Mux.scala 46:16:@12367.4]
  assign _T_15013 = 6'h24 == _T_10211_54; // @[Mux.scala 46:19:@12368.4]
  assign _T_15014 = _T_15013 ? _T_9260_35 : _T_15012; // @[Mux.scala 46:16:@12369.4]
  assign _T_15015 = 6'h23 == _T_10211_54; // @[Mux.scala 46:19:@12370.4]
  assign _T_15016 = _T_15015 ? _T_9260_34 : _T_15014; // @[Mux.scala 46:16:@12371.4]
  assign _T_15017 = 6'h22 == _T_10211_54; // @[Mux.scala 46:19:@12372.4]
  assign _T_15018 = _T_15017 ? _T_9260_33 : _T_15016; // @[Mux.scala 46:16:@12373.4]
  assign _T_15019 = 6'h21 == _T_10211_54; // @[Mux.scala 46:19:@12374.4]
  assign _T_15020 = _T_15019 ? _T_9260_32 : _T_15018; // @[Mux.scala 46:16:@12375.4]
  assign _T_15021 = 6'h20 == _T_10211_54; // @[Mux.scala 46:19:@12376.4]
  assign _T_15022 = _T_15021 ? _T_9260_31 : _T_15020; // @[Mux.scala 46:16:@12377.4]
  assign _T_15023 = 6'h1f == _T_10211_54; // @[Mux.scala 46:19:@12378.4]
  assign _T_15024 = _T_15023 ? _T_9260_30 : _T_15022; // @[Mux.scala 46:16:@12379.4]
  assign _T_15025 = 6'h1e == _T_10211_54; // @[Mux.scala 46:19:@12380.4]
  assign _T_15026 = _T_15025 ? _T_9260_29 : _T_15024; // @[Mux.scala 46:16:@12381.4]
  assign _T_15027 = 6'h1d == _T_10211_54; // @[Mux.scala 46:19:@12382.4]
  assign _T_15028 = _T_15027 ? _T_9260_28 : _T_15026; // @[Mux.scala 46:16:@12383.4]
  assign _T_15029 = 6'h1c == _T_10211_54; // @[Mux.scala 46:19:@12384.4]
  assign _T_15030 = _T_15029 ? _T_9260_27 : _T_15028; // @[Mux.scala 46:16:@12385.4]
  assign _T_15031 = 6'h1b == _T_10211_54; // @[Mux.scala 46:19:@12386.4]
  assign _T_15032 = _T_15031 ? _T_9260_26 : _T_15030; // @[Mux.scala 46:16:@12387.4]
  assign _T_15033 = 6'h1a == _T_10211_54; // @[Mux.scala 46:19:@12388.4]
  assign _T_15034 = _T_15033 ? _T_9260_25 : _T_15032; // @[Mux.scala 46:16:@12389.4]
  assign _T_15035 = 6'h19 == _T_10211_54; // @[Mux.scala 46:19:@12390.4]
  assign _T_15036 = _T_15035 ? _T_9260_24 : _T_15034; // @[Mux.scala 46:16:@12391.4]
  assign _T_15037 = 6'h18 == _T_10211_54; // @[Mux.scala 46:19:@12392.4]
  assign _T_15038 = _T_15037 ? _T_9260_23 : _T_15036; // @[Mux.scala 46:16:@12393.4]
  assign _T_15039 = 6'h17 == _T_10211_54; // @[Mux.scala 46:19:@12394.4]
  assign _T_15040 = _T_15039 ? _T_9260_22 : _T_15038; // @[Mux.scala 46:16:@12395.4]
  assign _T_15041 = 6'h16 == _T_10211_54; // @[Mux.scala 46:19:@12396.4]
  assign _T_15042 = _T_15041 ? _T_9260_21 : _T_15040; // @[Mux.scala 46:16:@12397.4]
  assign _T_15043 = 6'h15 == _T_10211_54; // @[Mux.scala 46:19:@12398.4]
  assign _T_15044 = _T_15043 ? _T_9260_20 : _T_15042; // @[Mux.scala 46:16:@12399.4]
  assign _T_15045 = 6'h14 == _T_10211_54; // @[Mux.scala 46:19:@12400.4]
  assign _T_15046 = _T_15045 ? _T_9260_19 : _T_15044; // @[Mux.scala 46:16:@12401.4]
  assign _T_15047 = 6'h13 == _T_10211_54; // @[Mux.scala 46:19:@12402.4]
  assign _T_15048 = _T_15047 ? _T_9260_18 : _T_15046; // @[Mux.scala 46:16:@12403.4]
  assign _T_15049 = 6'h12 == _T_10211_54; // @[Mux.scala 46:19:@12404.4]
  assign _T_15050 = _T_15049 ? _T_9260_17 : _T_15048; // @[Mux.scala 46:16:@12405.4]
  assign _T_15051 = 6'h11 == _T_10211_54; // @[Mux.scala 46:19:@12406.4]
  assign _T_15052 = _T_15051 ? _T_9260_16 : _T_15050; // @[Mux.scala 46:16:@12407.4]
  assign _T_15053 = 6'h10 == _T_10211_54; // @[Mux.scala 46:19:@12408.4]
  assign _T_15054 = _T_15053 ? _T_9260_15 : _T_15052; // @[Mux.scala 46:16:@12409.4]
  assign _T_15055 = 6'hf == _T_10211_54; // @[Mux.scala 46:19:@12410.4]
  assign _T_15056 = _T_15055 ? _T_9260_14 : _T_15054; // @[Mux.scala 46:16:@12411.4]
  assign _T_15057 = 6'he == _T_10211_54; // @[Mux.scala 46:19:@12412.4]
  assign _T_15058 = _T_15057 ? _T_9260_13 : _T_15056; // @[Mux.scala 46:16:@12413.4]
  assign _T_15059 = 6'hd == _T_10211_54; // @[Mux.scala 46:19:@12414.4]
  assign _T_15060 = _T_15059 ? _T_9260_12 : _T_15058; // @[Mux.scala 46:16:@12415.4]
  assign _T_15061 = 6'hc == _T_10211_54; // @[Mux.scala 46:19:@12416.4]
  assign _T_15062 = _T_15061 ? _T_9260_11 : _T_15060; // @[Mux.scala 46:16:@12417.4]
  assign _T_15063 = 6'hb == _T_10211_54; // @[Mux.scala 46:19:@12418.4]
  assign _T_15064 = _T_15063 ? _T_9260_10 : _T_15062; // @[Mux.scala 46:16:@12419.4]
  assign _T_15065 = 6'ha == _T_10211_54; // @[Mux.scala 46:19:@12420.4]
  assign _T_15066 = _T_15065 ? _T_9260_9 : _T_15064; // @[Mux.scala 46:16:@12421.4]
  assign _T_15067 = 6'h9 == _T_10211_54; // @[Mux.scala 46:19:@12422.4]
  assign _T_15068 = _T_15067 ? _T_9260_8 : _T_15066; // @[Mux.scala 46:16:@12423.4]
  assign _T_15069 = 6'h8 == _T_10211_54; // @[Mux.scala 46:19:@12424.4]
  assign _T_15070 = _T_15069 ? _T_9260_7 : _T_15068; // @[Mux.scala 46:16:@12425.4]
  assign _T_15071 = 6'h7 == _T_10211_54; // @[Mux.scala 46:19:@12426.4]
  assign _T_15072 = _T_15071 ? _T_9260_6 : _T_15070; // @[Mux.scala 46:16:@12427.4]
  assign _T_15073 = 6'h6 == _T_10211_54; // @[Mux.scala 46:19:@12428.4]
  assign _T_15074 = _T_15073 ? _T_9260_5 : _T_15072; // @[Mux.scala 46:16:@12429.4]
  assign _T_15075 = 6'h5 == _T_10211_54; // @[Mux.scala 46:19:@12430.4]
  assign _T_15076 = _T_15075 ? _T_9260_4 : _T_15074; // @[Mux.scala 46:16:@12431.4]
  assign _T_15077 = 6'h4 == _T_10211_54; // @[Mux.scala 46:19:@12432.4]
  assign _T_15078 = _T_15077 ? _T_9260_3 : _T_15076; // @[Mux.scala 46:16:@12433.4]
  assign _T_15079 = 6'h3 == _T_10211_54; // @[Mux.scala 46:19:@12434.4]
  assign _T_15080 = _T_15079 ? _T_9260_2 : _T_15078; // @[Mux.scala 46:16:@12435.4]
  assign _T_15081 = 6'h2 == _T_10211_54; // @[Mux.scala 46:19:@12436.4]
  assign _T_15082 = _T_15081 ? _T_9260_1 : _T_15080; // @[Mux.scala 46:16:@12437.4]
  assign _T_15083 = 6'h1 == _T_10211_54; // @[Mux.scala 46:19:@12438.4]
  assign _T_15084 = _T_15083 ? _T_9260_0 : _T_15082; // @[Mux.scala 46:16:@12439.4]
  assign _T_15142 = 6'h38 == _T_10211_55; // @[Mux.scala 46:19:@12441.4]
  assign _T_15143 = _T_15142 ? _T_9260_55 : 8'h0; // @[Mux.scala 46:16:@12442.4]
  assign _T_15144 = 6'h37 == _T_10211_55; // @[Mux.scala 46:19:@12443.4]
  assign _T_15145 = _T_15144 ? _T_9260_54 : _T_15143; // @[Mux.scala 46:16:@12444.4]
  assign _T_15146 = 6'h36 == _T_10211_55; // @[Mux.scala 46:19:@12445.4]
  assign _T_15147 = _T_15146 ? _T_9260_53 : _T_15145; // @[Mux.scala 46:16:@12446.4]
  assign _T_15148 = 6'h35 == _T_10211_55; // @[Mux.scala 46:19:@12447.4]
  assign _T_15149 = _T_15148 ? _T_9260_52 : _T_15147; // @[Mux.scala 46:16:@12448.4]
  assign _T_15150 = 6'h34 == _T_10211_55; // @[Mux.scala 46:19:@12449.4]
  assign _T_15151 = _T_15150 ? _T_9260_51 : _T_15149; // @[Mux.scala 46:16:@12450.4]
  assign _T_15152 = 6'h33 == _T_10211_55; // @[Mux.scala 46:19:@12451.4]
  assign _T_15153 = _T_15152 ? _T_9260_50 : _T_15151; // @[Mux.scala 46:16:@12452.4]
  assign _T_15154 = 6'h32 == _T_10211_55; // @[Mux.scala 46:19:@12453.4]
  assign _T_15155 = _T_15154 ? _T_9260_49 : _T_15153; // @[Mux.scala 46:16:@12454.4]
  assign _T_15156 = 6'h31 == _T_10211_55; // @[Mux.scala 46:19:@12455.4]
  assign _T_15157 = _T_15156 ? _T_9260_48 : _T_15155; // @[Mux.scala 46:16:@12456.4]
  assign _T_15158 = 6'h30 == _T_10211_55; // @[Mux.scala 46:19:@12457.4]
  assign _T_15159 = _T_15158 ? _T_9260_47 : _T_15157; // @[Mux.scala 46:16:@12458.4]
  assign _T_15160 = 6'h2f == _T_10211_55; // @[Mux.scala 46:19:@12459.4]
  assign _T_15161 = _T_15160 ? _T_9260_46 : _T_15159; // @[Mux.scala 46:16:@12460.4]
  assign _T_15162 = 6'h2e == _T_10211_55; // @[Mux.scala 46:19:@12461.4]
  assign _T_15163 = _T_15162 ? _T_9260_45 : _T_15161; // @[Mux.scala 46:16:@12462.4]
  assign _T_15164 = 6'h2d == _T_10211_55; // @[Mux.scala 46:19:@12463.4]
  assign _T_15165 = _T_15164 ? _T_9260_44 : _T_15163; // @[Mux.scala 46:16:@12464.4]
  assign _T_15166 = 6'h2c == _T_10211_55; // @[Mux.scala 46:19:@12465.4]
  assign _T_15167 = _T_15166 ? _T_9260_43 : _T_15165; // @[Mux.scala 46:16:@12466.4]
  assign _T_15168 = 6'h2b == _T_10211_55; // @[Mux.scala 46:19:@12467.4]
  assign _T_15169 = _T_15168 ? _T_9260_42 : _T_15167; // @[Mux.scala 46:16:@12468.4]
  assign _T_15170 = 6'h2a == _T_10211_55; // @[Mux.scala 46:19:@12469.4]
  assign _T_15171 = _T_15170 ? _T_9260_41 : _T_15169; // @[Mux.scala 46:16:@12470.4]
  assign _T_15172 = 6'h29 == _T_10211_55; // @[Mux.scala 46:19:@12471.4]
  assign _T_15173 = _T_15172 ? _T_9260_40 : _T_15171; // @[Mux.scala 46:16:@12472.4]
  assign _T_15174 = 6'h28 == _T_10211_55; // @[Mux.scala 46:19:@12473.4]
  assign _T_15175 = _T_15174 ? _T_9260_39 : _T_15173; // @[Mux.scala 46:16:@12474.4]
  assign _T_15176 = 6'h27 == _T_10211_55; // @[Mux.scala 46:19:@12475.4]
  assign _T_15177 = _T_15176 ? _T_9260_38 : _T_15175; // @[Mux.scala 46:16:@12476.4]
  assign _T_15178 = 6'h26 == _T_10211_55; // @[Mux.scala 46:19:@12477.4]
  assign _T_15179 = _T_15178 ? _T_9260_37 : _T_15177; // @[Mux.scala 46:16:@12478.4]
  assign _T_15180 = 6'h25 == _T_10211_55; // @[Mux.scala 46:19:@12479.4]
  assign _T_15181 = _T_15180 ? _T_9260_36 : _T_15179; // @[Mux.scala 46:16:@12480.4]
  assign _T_15182 = 6'h24 == _T_10211_55; // @[Mux.scala 46:19:@12481.4]
  assign _T_15183 = _T_15182 ? _T_9260_35 : _T_15181; // @[Mux.scala 46:16:@12482.4]
  assign _T_15184 = 6'h23 == _T_10211_55; // @[Mux.scala 46:19:@12483.4]
  assign _T_15185 = _T_15184 ? _T_9260_34 : _T_15183; // @[Mux.scala 46:16:@12484.4]
  assign _T_15186 = 6'h22 == _T_10211_55; // @[Mux.scala 46:19:@12485.4]
  assign _T_15187 = _T_15186 ? _T_9260_33 : _T_15185; // @[Mux.scala 46:16:@12486.4]
  assign _T_15188 = 6'h21 == _T_10211_55; // @[Mux.scala 46:19:@12487.4]
  assign _T_15189 = _T_15188 ? _T_9260_32 : _T_15187; // @[Mux.scala 46:16:@12488.4]
  assign _T_15190 = 6'h20 == _T_10211_55; // @[Mux.scala 46:19:@12489.4]
  assign _T_15191 = _T_15190 ? _T_9260_31 : _T_15189; // @[Mux.scala 46:16:@12490.4]
  assign _T_15192 = 6'h1f == _T_10211_55; // @[Mux.scala 46:19:@12491.4]
  assign _T_15193 = _T_15192 ? _T_9260_30 : _T_15191; // @[Mux.scala 46:16:@12492.4]
  assign _T_15194 = 6'h1e == _T_10211_55; // @[Mux.scala 46:19:@12493.4]
  assign _T_15195 = _T_15194 ? _T_9260_29 : _T_15193; // @[Mux.scala 46:16:@12494.4]
  assign _T_15196 = 6'h1d == _T_10211_55; // @[Mux.scala 46:19:@12495.4]
  assign _T_15197 = _T_15196 ? _T_9260_28 : _T_15195; // @[Mux.scala 46:16:@12496.4]
  assign _T_15198 = 6'h1c == _T_10211_55; // @[Mux.scala 46:19:@12497.4]
  assign _T_15199 = _T_15198 ? _T_9260_27 : _T_15197; // @[Mux.scala 46:16:@12498.4]
  assign _T_15200 = 6'h1b == _T_10211_55; // @[Mux.scala 46:19:@12499.4]
  assign _T_15201 = _T_15200 ? _T_9260_26 : _T_15199; // @[Mux.scala 46:16:@12500.4]
  assign _T_15202 = 6'h1a == _T_10211_55; // @[Mux.scala 46:19:@12501.4]
  assign _T_15203 = _T_15202 ? _T_9260_25 : _T_15201; // @[Mux.scala 46:16:@12502.4]
  assign _T_15204 = 6'h19 == _T_10211_55; // @[Mux.scala 46:19:@12503.4]
  assign _T_15205 = _T_15204 ? _T_9260_24 : _T_15203; // @[Mux.scala 46:16:@12504.4]
  assign _T_15206 = 6'h18 == _T_10211_55; // @[Mux.scala 46:19:@12505.4]
  assign _T_15207 = _T_15206 ? _T_9260_23 : _T_15205; // @[Mux.scala 46:16:@12506.4]
  assign _T_15208 = 6'h17 == _T_10211_55; // @[Mux.scala 46:19:@12507.4]
  assign _T_15209 = _T_15208 ? _T_9260_22 : _T_15207; // @[Mux.scala 46:16:@12508.4]
  assign _T_15210 = 6'h16 == _T_10211_55; // @[Mux.scala 46:19:@12509.4]
  assign _T_15211 = _T_15210 ? _T_9260_21 : _T_15209; // @[Mux.scala 46:16:@12510.4]
  assign _T_15212 = 6'h15 == _T_10211_55; // @[Mux.scala 46:19:@12511.4]
  assign _T_15213 = _T_15212 ? _T_9260_20 : _T_15211; // @[Mux.scala 46:16:@12512.4]
  assign _T_15214 = 6'h14 == _T_10211_55; // @[Mux.scala 46:19:@12513.4]
  assign _T_15215 = _T_15214 ? _T_9260_19 : _T_15213; // @[Mux.scala 46:16:@12514.4]
  assign _T_15216 = 6'h13 == _T_10211_55; // @[Mux.scala 46:19:@12515.4]
  assign _T_15217 = _T_15216 ? _T_9260_18 : _T_15215; // @[Mux.scala 46:16:@12516.4]
  assign _T_15218 = 6'h12 == _T_10211_55; // @[Mux.scala 46:19:@12517.4]
  assign _T_15219 = _T_15218 ? _T_9260_17 : _T_15217; // @[Mux.scala 46:16:@12518.4]
  assign _T_15220 = 6'h11 == _T_10211_55; // @[Mux.scala 46:19:@12519.4]
  assign _T_15221 = _T_15220 ? _T_9260_16 : _T_15219; // @[Mux.scala 46:16:@12520.4]
  assign _T_15222 = 6'h10 == _T_10211_55; // @[Mux.scala 46:19:@12521.4]
  assign _T_15223 = _T_15222 ? _T_9260_15 : _T_15221; // @[Mux.scala 46:16:@12522.4]
  assign _T_15224 = 6'hf == _T_10211_55; // @[Mux.scala 46:19:@12523.4]
  assign _T_15225 = _T_15224 ? _T_9260_14 : _T_15223; // @[Mux.scala 46:16:@12524.4]
  assign _T_15226 = 6'he == _T_10211_55; // @[Mux.scala 46:19:@12525.4]
  assign _T_15227 = _T_15226 ? _T_9260_13 : _T_15225; // @[Mux.scala 46:16:@12526.4]
  assign _T_15228 = 6'hd == _T_10211_55; // @[Mux.scala 46:19:@12527.4]
  assign _T_15229 = _T_15228 ? _T_9260_12 : _T_15227; // @[Mux.scala 46:16:@12528.4]
  assign _T_15230 = 6'hc == _T_10211_55; // @[Mux.scala 46:19:@12529.4]
  assign _T_15231 = _T_15230 ? _T_9260_11 : _T_15229; // @[Mux.scala 46:16:@12530.4]
  assign _T_15232 = 6'hb == _T_10211_55; // @[Mux.scala 46:19:@12531.4]
  assign _T_15233 = _T_15232 ? _T_9260_10 : _T_15231; // @[Mux.scala 46:16:@12532.4]
  assign _T_15234 = 6'ha == _T_10211_55; // @[Mux.scala 46:19:@12533.4]
  assign _T_15235 = _T_15234 ? _T_9260_9 : _T_15233; // @[Mux.scala 46:16:@12534.4]
  assign _T_15236 = 6'h9 == _T_10211_55; // @[Mux.scala 46:19:@12535.4]
  assign _T_15237 = _T_15236 ? _T_9260_8 : _T_15235; // @[Mux.scala 46:16:@12536.4]
  assign _T_15238 = 6'h8 == _T_10211_55; // @[Mux.scala 46:19:@12537.4]
  assign _T_15239 = _T_15238 ? _T_9260_7 : _T_15237; // @[Mux.scala 46:16:@12538.4]
  assign _T_15240 = 6'h7 == _T_10211_55; // @[Mux.scala 46:19:@12539.4]
  assign _T_15241 = _T_15240 ? _T_9260_6 : _T_15239; // @[Mux.scala 46:16:@12540.4]
  assign _T_15242 = 6'h6 == _T_10211_55; // @[Mux.scala 46:19:@12541.4]
  assign _T_15243 = _T_15242 ? _T_9260_5 : _T_15241; // @[Mux.scala 46:16:@12542.4]
  assign _T_15244 = 6'h5 == _T_10211_55; // @[Mux.scala 46:19:@12543.4]
  assign _T_15245 = _T_15244 ? _T_9260_4 : _T_15243; // @[Mux.scala 46:16:@12544.4]
  assign _T_15246 = 6'h4 == _T_10211_55; // @[Mux.scala 46:19:@12545.4]
  assign _T_15247 = _T_15246 ? _T_9260_3 : _T_15245; // @[Mux.scala 46:16:@12546.4]
  assign _T_15248 = 6'h3 == _T_10211_55; // @[Mux.scala 46:19:@12547.4]
  assign _T_15249 = _T_15248 ? _T_9260_2 : _T_15247; // @[Mux.scala 46:16:@12548.4]
  assign _T_15250 = 6'h2 == _T_10211_55; // @[Mux.scala 46:19:@12549.4]
  assign _T_15251 = _T_15250 ? _T_9260_1 : _T_15249; // @[Mux.scala 46:16:@12550.4]
  assign _T_15252 = 6'h1 == _T_10211_55; // @[Mux.scala 46:19:@12551.4]
  assign _T_15253 = _T_15252 ? _T_9260_0 : _T_15251; // @[Mux.scala 46:16:@12552.4]
  assign _T_15312 = 6'h39 == _T_10211_56; // @[Mux.scala 46:19:@12554.4]
  assign _T_15313 = _T_15312 ? _T_9260_56 : 8'h0; // @[Mux.scala 46:16:@12555.4]
  assign _T_15314 = 6'h38 == _T_10211_56; // @[Mux.scala 46:19:@12556.4]
  assign _T_15315 = _T_15314 ? _T_9260_55 : _T_15313; // @[Mux.scala 46:16:@12557.4]
  assign _T_15316 = 6'h37 == _T_10211_56; // @[Mux.scala 46:19:@12558.4]
  assign _T_15317 = _T_15316 ? _T_9260_54 : _T_15315; // @[Mux.scala 46:16:@12559.4]
  assign _T_15318 = 6'h36 == _T_10211_56; // @[Mux.scala 46:19:@12560.4]
  assign _T_15319 = _T_15318 ? _T_9260_53 : _T_15317; // @[Mux.scala 46:16:@12561.4]
  assign _T_15320 = 6'h35 == _T_10211_56; // @[Mux.scala 46:19:@12562.4]
  assign _T_15321 = _T_15320 ? _T_9260_52 : _T_15319; // @[Mux.scala 46:16:@12563.4]
  assign _T_15322 = 6'h34 == _T_10211_56; // @[Mux.scala 46:19:@12564.4]
  assign _T_15323 = _T_15322 ? _T_9260_51 : _T_15321; // @[Mux.scala 46:16:@12565.4]
  assign _T_15324 = 6'h33 == _T_10211_56; // @[Mux.scala 46:19:@12566.4]
  assign _T_15325 = _T_15324 ? _T_9260_50 : _T_15323; // @[Mux.scala 46:16:@12567.4]
  assign _T_15326 = 6'h32 == _T_10211_56; // @[Mux.scala 46:19:@12568.4]
  assign _T_15327 = _T_15326 ? _T_9260_49 : _T_15325; // @[Mux.scala 46:16:@12569.4]
  assign _T_15328 = 6'h31 == _T_10211_56; // @[Mux.scala 46:19:@12570.4]
  assign _T_15329 = _T_15328 ? _T_9260_48 : _T_15327; // @[Mux.scala 46:16:@12571.4]
  assign _T_15330 = 6'h30 == _T_10211_56; // @[Mux.scala 46:19:@12572.4]
  assign _T_15331 = _T_15330 ? _T_9260_47 : _T_15329; // @[Mux.scala 46:16:@12573.4]
  assign _T_15332 = 6'h2f == _T_10211_56; // @[Mux.scala 46:19:@12574.4]
  assign _T_15333 = _T_15332 ? _T_9260_46 : _T_15331; // @[Mux.scala 46:16:@12575.4]
  assign _T_15334 = 6'h2e == _T_10211_56; // @[Mux.scala 46:19:@12576.4]
  assign _T_15335 = _T_15334 ? _T_9260_45 : _T_15333; // @[Mux.scala 46:16:@12577.4]
  assign _T_15336 = 6'h2d == _T_10211_56; // @[Mux.scala 46:19:@12578.4]
  assign _T_15337 = _T_15336 ? _T_9260_44 : _T_15335; // @[Mux.scala 46:16:@12579.4]
  assign _T_15338 = 6'h2c == _T_10211_56; // @[Mux.scala 46:19:@12580.4]
  assign _T_15339 = _T_15338 ? _T_9260_43 : _T_15337; // @[Mux.scala 46:16:@12581.4]
  assign _T_15340 = 6'h2b == _T_10211_56; // @[Mux.scala 46:19:@12582.4]
  assign _T_15341 = _T_15340 ? _T_9260_42 : _T_15339; // @[Mux.scala 46:16:@12583.4]
  assign _T_15342 = 6'h2a == _T_10211_56; // @[Mux.scala 46:19:@12584.4]
  assign _T_15343 = _T_15342 ? _T_9260_41 : _T_15341; // @[Mux.scala 46:16:@12585.4]
  assign _T_15344 = 6'h29 == _T_10211_56; // @[Mux.scala 46:19:@12586.4]
  assign _T_15345 = _T_15344 ? _T_9260_40 : _T_15343; // @[Mux.scala 46:16:@12587.4]
  assign _T_15346 = 6'h28 == _T_10211_56; // @[Mux.scala 46:19:@12588.4]
  assign _T_15347 = _T_15346 ? _T_9260_39 : _T_15345; // @[Mux.scala 46:16:@12589.4]
  assign _T_15348 = 6'h27 == _T_10211_56; // @[Mux.scala 46:19:@12590.4]
  assign _T_15349 = _T_15348 ? _T_9260_38 : _T_15347; // @[Mux.scala 46:16:@12591.4]
  assign _T_15350 = 6'h26 == _T_10211_56; // @[Mux.scala 46:19:@12592.4]
  assign _T_15351 = _T_15350 ? _T_9260_37 : _T_15349; // @[Mux.scala 46:16:@12593.4]
  assign _T_15352 = 6'h25 == _T_10211_56; // @[Mux.scala 46:19:@12594.4]
  assign _T_15353 = _T_15352 ? _T_9260_36 : _T_15351; // @[Mux.scala 46:16:@12595.4]
  assign _T_15354 = 6'h24 == _T_10211_56; // @[Mux.scala 46:19:@12596.4]
  assign _T_15355 = _T_15354 ? _T_9260_35 : _T_15353; // @[Mux.scala 46:16:@12597.4]
  assign _T_15356 = 6'h23 == _T_10211_56; // @[Mux.scala 46:19:@12598.4]
  assign _T_15357 = _T_15356 ? _T_9260_34 : _T_15355; // @[Mux.scala 46:16:@12599.4]
  assign _T_15358 = 6'h22 == _T_10211_56; // @[Mux.scala 46:19:@12600.4]
  assign _T_15359 = _T_15358 ? _T_9260_33 : _T_15357; // @[Mux.scala 46:16:@12601.4]
  assign _T_15360 = 6'h21 == _T_10211_56; // @[Mux.scala 46:19:@12602.4]
  assign _T_15361 = _T_15360 ? _T_9260_32 : _T_15359; // @[Mux.scala 46:16:@12603.4]
  assign _T_15362 = 6'h20 == _T_10211_56; // @[Mux.scala 46:19:@12604.4]
  assign _T_15363 = _T_15362 ? _T_9260_31 : _T_15361; // @[Mux.scala 46:16:@12605.4]
  assign _T_15364 = 6'h1f == _T_10211_56; // @[Mux.scala 46:19:@12606.4]
  assign _T_15365 = _T_15364 ? _T_9260_30 : _T_15363; // @[Mux.scala 46:16:@12607.4]
  assign _T_15366 = 6'h1e == _T_10211_56; // @[Mux.scala 46:19:@12608.4]
  assign _T_15367 = _T_15366 ? _T_9260_29 : _T_15365; // @[Mux.scala 46:16:@12609.4]
  assign _T_15368 = 6'h1d == _T_10211_56; // @[Mux.scala 46:19:@12610.4]
  assign _T_15369 = _T_15368 ? _T_9260_28 : _T_15367; // @[Mux.scala 46:16:@12611.4]
  assign _T_15370 = 6'h1c == _T_10211_56; // @[Mux.scala 46:19:@12612.4]
  assign _T_15371 = _T_15370 ? _T_9260_27 : _T_15369; // @[Mux.scala 46:16:@12613.4]
  assign _T_15372 = 6'h1b == _T_10211_56; // @[Mux.scala 46:19:@12614.4]
  assign _T_15373 = _T_15372 ? _T_9260_26 : _T_15371; // @[Mux.scala 46:16:@12615.4]
  assign _T_15374 = 6'h1a == _T_10211_56; // @[Mux.scala 46:19:@12616.4]
  assign _T_15375 = _T_15374 ? _T_9260_25 : _T_15373; // @[Mux.scala 46:16:@12617.4]
  assign _T_15376 = 6'h19 == _T_10211_56; // @[Mux.scala 46:19:@12618.4]
  assign _T_15377 = _T_15376 ? _T_9260_24 : _T_15375; // @[Mux.scala 46:16:@12619.4]
  assign _T_15378 = 6'h18 == _T_10211_56; // @[Mux.scala 46:19:@12620.4]
  assign _T_15379 = _T_15378 ? _T_9260_23 : _T_15377; // @[Mux.scala 46:16:@12621.4]
  assign _T_15380 = 6'h17 == _T_10211_56; // @[Mux.scala 46:19:@12622.4]
  assign _T_15381 = _T_15380 ? _T_9260_22 : _T_15379; // @[Mux.scala 46:16:@12623.4]
  assign _T_15382 = 6'h16 == _T_10211_56; // @[Mux.scala 46:19:@12624.4]
  assign _T_15383 = _T_15382 ? _T_9260_21 : _T_15381; // @[Mux.scala 46:16:@12625.4]
  assign _T_15384 = 6'h15 == _T_10211_56; // @[Mux.scala 46:19:@12626.4]
  assign _T_15385 = _T_15384 ? _T_9260_20 : _T_15383; // @[Mux.scala 46:16:@12627.4]
  assign _T_15386 = 6'h14 == _T_10211_56; // @[Mux.scala 46:19:@12628.4]
  assign _T_15387 = _T_15386 ? _T_9260_19 : _T_15385; // @[Mux.scala 46:16:@12629.4]
  assign _T_15388 = 6'h13 == _T_10211_56; // @[Mux.scala 46:19:@12630.4]
  assign _T_15389 = _T_15388 ? _T_9260_18 : _T_15387; // @[Mux.scala 46:16:@12631.4]
  assign _T_15390 = 6'h12 == _T_10211_56; // @[Mux.scala 46:19:@12632.4]
  assign _T_15391 = _T_15390 ? _T_9260_17 : _T_15389; // @[Mux.scala 46:16:@12633.4]
  assign _T_15392 = 6'h11 == _T_10211_56; // @[Mux.scala 46:19:@12634.4]
  assign _T_15393 = _T_15392 ? _T_9260_16 : _T_15391; // @[Mux.scala 46:16:@12635.4]
  assign _T_15394 = 6'h10 == _T_10211_56; // @[Mux.scala 46:19:@12636.4]
  assign _T_15395 = _T_15394 ? _T_9260_15 : _T_15393; // @[Mux.scala 46:16:@12637.4]
  assign _T_15396 = 6'hf == _T_10211_56; // @[Mux.scala 46:19:@12638.4]
  assign _T_15397 = _T_15396 ? _T_9260_14 : _T_15395; // @[Mux.scala 46:16:@12639.4]
  assign _T_15398 = 6'he == _T_10211_56; // @[Mux.scala 46:19:@12640.4]
  assign _T_15399 = _T_15398 ? _T_9260_13 : _T_15397; // @[Mux.scala 46:16:@12641.4]
  assign _T_15400 = 6'hd == _T_10211_56; // @[Mux.scala 46:19:@12642.4]
  assign _T_15401 = _T_15400 ? _T_9260_12 : _T_15399; // @[Mux.scala 46:16:@12643.4]
  assign _T_15402 = 6'hc == _T_10211_56; // @[Mux.scala 46:19:@12644.4]
  assign _T_15403 = _T_15402 ? _T_9260_11 : _T_15401; // @[Mux.scala 46:16:@12645.4]
  assign _T_15404 = 6'hb == _T_10211_56; // @[Mux.scala 46:19:@12646.4]
  assign _T_15405 = _T_15404 ? _T_9260_10 : _T_15403; // @[Mux.scala 46:16:@12647.4]
  assign _T_15406 = 6'ha == _T_10211_56; // @[Mux.scala 46:19:@12648.4]
  assign _T_15407 = _T_15406 ? _T_9260_9 : _T_15405; // @[Mux.scala 46:16:@12649.4]
  assign _T_15408 = 6'h9 == _T_10211_56; // @[Mux.scala 46:19:@12650.4]
  assign _T_15409 = _T_15408 ? _T_9260_8 : _T_15407; // @[Mux.scala 46:16:@12651.4]
  assign _T_15410 = 6'h8 == _T_10211_56; // @[Mux.scala 46:19:@12652.4]
  assign _T_15411 = _T_15410 ? _T_9260_7 : _T_15409; // @[Mux.scala 46:16:@12653.4]
  assign _T_15412 = 6'h7 == _T_10211_56; // @[Mux.scala 46:19:@12654.4]
  assign _T_15413 = _T_15412 ? _T_9260_6 : _T_15411; // @[Mux.scala 46:16:@12655.4]
  assign _T_15414 = 6'h6 == _T_10211_56; // @[Mux.scala 46:19:@12656.4]
  assign _T_15415 = _T_15414 ? _T_9260_5 : _T_15413; // @[Mux.scala 46:16:@12657.4]
  assign _T_15416 = 6'h5 == _T_10211_56; // @[Mux.scala 46:19:@12658.4]
  assign _T_15417 = _T_15416 ? _T_9260_4 : _T_15415; // @[Mux.scala 46:16:@12659.4]
  assign _T_15418 = 6'h4 == _T_10211_56; // @[Mux.scala 46:19:@12660.4]
  assign _T_15419 = _T_15418 ? _T_9260_3 : _T_15417; // @[Mux.scala 46:16:@12661.4]
  assign _T_15420 = 6'h3 == _T_10211_56; // @[Mux.scala 46:19:@12662.4]
  assign _T_15421 = _T_15420 ? _T_9260_2 : _T_15419; // @[Mux.scala 46:16:@12663.4]
  assign _T_15422 = 6'h2 == _T_10211_56; // @[Mux.scala 46:19:@12664.4]
  assign _T_15423 = _T_15422 ? _T_9260_1 : _T_15421; // @[Mux.scala 46:16:@12665.4]
  assign _T_15424 = 6'h1 == _T_10211_56; // @[Mux.scala 46:19:@12666.4]
  assign _T_15425 = _T_15424 ? _T_9260_0 : _T_15423; // @[Mux.scala 46:16:@12667.4]
  assign _T_15485 = 6'h3a == _T_10211_57; // @[Mux.scala 46:19:@12669.4]
  assign _T_15486 = _T_15485 ? _T_9260_57 : 8'h0; // @[Mux.scala 46:16:@12670.4]
  assign _T_15487 = 6'h39 == _T_10211_57; // @[Mux.scala 46:19:@12671.4]
  assign _T_15488 = _T_15487 ? _T_9260_56 : _T_15486; // @[Mux.scala 46:16:@12672.4]
  assign _T_15489 = 6'h38 == _T_10211_57; // @[Mux.scala 46:19:@12673.4]
  assign _T_15490 = _T_15489 ? _T_9260_55 : _T_15488; // @[Mux.scala 46:16:@12674.4]
  assign _T_15491 = 6'h37 == _T_10211_57; // @[Mux.scala 46:19:@12675.4]
  assign _T_15492 = _T_15491 ? _T_9260_54 : _T_15490; // @[Mux.scala 46:16:@12676.4]
  assign _T_15493 = 6'h36 == _T_10211_57; // @[Mux.scala 46:19:@12677.4]
  assign _T_15494 = _T_15493 ? _T_9260_53 : _T_15492; // @[Mux.scala 46:16:@12678.4]
  assign _T_15495 = 6'h35 == _T_10211_57; // @[Mux.scala 46:19:@12679.4]
  assign _T_15496 = _T_15495 ? _T_9260_52 : _T_15494; // @[Mux.scala 46:16:@12680.4]
  assign _T_15497 = 6'h34 == _T_10211_57; // @[Mux.scala 46:19:@12681.4]
  assign _T_15498 = _T_15497 ? _T_9260_51 : _T_15496; // @[Mux.scala 46:16:@12682.4]
  assign _T_15499 = 6'h33 == _T_10211_57; // @[Mux.scala 46:19:@12683.4]
  assign _T_15500 = _T_15499 ? _T_9260_50 : _T_15498; // @[Mux.scala 46:16:@12684.4]
  assign _T_15501 = 6'h32 == _T_10211_57; // @[Mux.scala 46:19:@12685.4]
  assign _T_15502 = _T_15501 ? _T_9260_49 : _T_15500; // @[Mux.scala 46:16:@12686.4]
  assign _T_15503 = 6'h31 == _T_10211_57; // @[Mux.scala 46:19:@12687.4]
  assign _T_15504 = _T_15503 ? _T_9260_48 : _T_15502; // @[Mux.scala 46:16:@12688.4]
  assign _T_15505 = 6'h30 == _T_10211_57; // @[Mux.scala 46:19:@12689.4]
  assign _T_15506 = _T_15505 ? _T_9260_47 : _T_15504; // @[Mux.scala 46:16:@12690.4]
  assign _T_15507 = 6'h2f == _T_10211_57; // @[Mux.scala 46:19:@12691.4]
  assign _T_15508 = _T_15507 ? _T_9260_46 : _T_15506; // @[Mux.scala 46:16:@12692.4]
  assign _T_15509 = 6'h2e == _T_10211_57; // @[Mux.scala 46:19:@12693.4]
  assign _T_15510 = _T_15509 ? _T_9260_45 : _T_15508; // @[Mux.scala 46:16:@12694.4]
  assign _T_15511 = 6'h2d == _T_10211_57; // @[Mux.scala 46:19:@12695.4]
  assign _T_15512 = _T_15511 ? _T_9260_44 : _T_15510; // @[Mux.scala 46:16:@12696.4]
  assign _T_15513 = 6'h2c == _T_10211_57; // @[Mux.scala 46:19:@12697.4]
  assign _T_15514 = _T_15513 ? _T_9260_43 : _T_15512; // @[Mux.scala 46:16:@12698.4]
  assign _T_15515 = 6'h2b == _T_10211_57; // @[Mux.scala 46:19:@12699.4]
  assign _T_15516 = _T_15515 ? _T_9260_42 : _T_15514; // @[Mux.scala 46:16:@12700.4]
  assign _T_15517 = 6'h2a == _T_10211_57; // @[Mux.scala 46:19:@12701.4]
  assign _T_15518 = _T_15517 ? _T_9260_41 : _T_15516; // @[Mux.scala 46:16:@12702.4]
  assign _T_15519 = 6'h29 == _T_10211_57; // @[Mux.scala 46:19:@12703.4]
  assign _T_15520 = _T_15519 ? _T_9260_40 : _T_15518; // @[Mux.scala 46:16:@12704.4]
  assign _T_15521 = 6'h28 == _T_10211_57; // @[Mux.scala 46:19:@12705.4]
  assign _T_15522 = _T_15521 ? _T_9260_39 : _T_15520; // @[Mux.scala 46:16:@12706.4]
  assign _T_15523 = 6'h27 == _T_10211_57; // @[Mux.scala 46:19:@12707.4]
  assign _T_15524 = _T_15523 ? _T_9260_38 : _T_15522; // @[Mux.scala 46:16:@12708.4]
  assign _T_15525 = 6'h26 == _T_10211_57; // @[Mux.scala 46:19:@12709.4]
  assign _T_15526 = _T_15525 ? _T_9260_37 : _T_15524; // @[Mux.scala 46:16:@12710.4]
  assign _T_15527 = 6'h25 == _T_10211_57; // @[Mux.scala 46:19:@12711.4]
  assign _T_15528 = _T_15527 ? _T_9260_36 : _T_15526; // @[Mux.scala 46:16:@12712.4]
  assign _T_15529 = 6'h24 == _T_10211_57; // @[Mux.scala 46:19:@12713.4]
  assign _T_15530 = _T_15529 ? _T_9260_35 : _T_15528; // @[Mux.scala 46:16:@12714.4]
  assign _T_15531 = 6'h23 == _T_10211_57; // @[Mux.scala 46:19:@12715.4]
  assign _T_15532 = _T_15531 ? _T_9260_34 : _T_15530; // @[Mux.scala 46:16:@12716.4]
  assign _T_15533 = 6'h22 == _T_10211_57; // @[Mux.scala 46:19:@12717.4]
  assign _T_15534 = _T_15533 ? _T_9260_33 : _T_15532; // @[Mux.scala 46:16:@12718.4]
  assign _T_15535 = 6'h21 == _T_10211_57; // @[Mux.scala 46:19:@12719.4]
  assign _T_15536 = _T_15535 ? _T_9260_32 : _T_15534; // @[Mux.scala 46:16:@12720.4]
  assign _T_15537 = 6'h20 == _T_10211_57; // @[Mux.scala 46:19:@12721.4]
  assign _T_15538 = _T_15537 ? _T_9260_31 : _T_15536; // @[Mux.scala 46:16:@12722.4]
  assign _T_15539 = 6'h1f == _T_10211_57; // @[Mux.scala 46:19:@12723.4]
  assign _T_15540 = _T_15539 ? _T_9260_30 : _T_15538; // @[Mux.scala 46:16:@12724.4]
  assign _T_15541 = 6'h1e == _T_10211_57; // @[Mux.scala 46:19:@12725.4]
  assign _T_15542 = _T_15541 ? _T_9260_29 : _T_15540; // @[Mux.scala 46:16:@12726.4]
  assign _T_15543 = 6'h1d == _T_10211_57; // @[Mux.scala 46:19:@12727.4]
  assign _T_15544 = _T_15543 ? _T_9260_28 : _T_15542; // @[Mux.scala 46:16:@12728.4]
  assign _T_15545 = 6'h1c == _T_10211_57; // @[Mux.scala 46:19:@12729.4]
  assign _T_15546 = _T_15545 ? _T_9260_27 : _T_15544; // @[Mux.scala 46:16:@12730.4]
  assign _T_15547 = 6'h1b == _T_10211_57; // @[Mux.scala 46:19:@12731.4]
  assign _T_15548 = _T_15547 ? _T_9260_26 : _T_15546; // @[Mux.scala 46:16:@12732.4]
  assign _T_15549 = 6'h1a == _T_10211_57; // @[Mux.scala 46:19:@12733.4]
  assign _T_15550 = _T_15549 ? _T_9260_25 : _T_15548; // @[Mux.scala 46:16:@12734.4]
  assign _T_15551 = 6'h19 == _T_10211_57; // @[Mux.scala 46:19:@12735.4]
  assign _T_15552 = _T_15551 ? _T_9260_24 : _T_15550; // @[Mux.scala 46:16:@12736.4]
  assign _T_15553 = 6'h18 == _T_10211_57; // @[Mux.scala 46:19:@12737.4]
  assign _T_15554 = _T_15553 ? _T_9260_23 : _T_15552; // @[Mux.scala 46:16:@12738.4]
  assign _T_15555 = 6'h17 == _T_10211_57; // @[Mux.scala 46:19:@12739.4]
  assign _T_15556 = _T_15555 ? _T_9260_22 : _T_15554; // @[Mux.scala 46:16:@12740.4]
  assign _T_15557 = 6'h16 == _T_10211_57; // @[Mux.scala 46:19:@12741.4]
  assign _T_15558 = _T_15557 ? _T_9260_21 : _T_15556; // @[Mux.scala 46:16:@12742.4]
  assign _T_15559 = 6'h15 == _T_10211_57; // @[Mux.scala 46:19:@12743.4]
  assign _T_15560 = _T_15559 ? _T_9260_20 : _T_15558; // @[Mux.scala 46:16:@12744.4]
  assign _T_15561 = 6'h14 == _T_10211_57; // @[Mux.scala 46:19:@12745.4]
  assign _T_15562 = _T_15561 ? _T_9260_19 : _T_15560; // @[Mux.scala 46:16:@12746.4]
  assign _T_15563 = 6'h13 == _T_10211_57; // @[Mux.scala 46:19:@12747.4]
  assign _T_15564 = _T_15563 ? _T_9260_18 : _T_15562; // @[Mux.scala 46:16:@12748.4]
  assign _T_15565 = 6'h12 == _T_10211_57; // @[Mux.scala 46:19:@12749.4]
  assign _T_15566 = _T_15565 ? _T_9260_17 : _T_15564; // @[Mux.scala 46:16:@12750.4]
  assign _T_15567 = 6'h11 == _T_10211_57; // @[Mux.scala 46:19:@12751.4]
  assign _T_15568 = _T_15567 ? _T_9260_16 : _T_15566; // @[Mux.scala 46:16:@12752.4]
  assign _T_15569 = 6'h10 == _T_10211_57; // @[Mux.scala 46:19:@12753.4]
  assign _T_15570 = _T_15569 ? _T_9260_15 : _T_15568; // @[Mux.scala 46:16:@12754.4]
  assign _T_15571 = 6'hf == _T_10211_57; // @[Mux.scala 46:19:@12755.4]
  assign _T_15572 = _T_15571 ? _T_9260_14 : _T_15570; // @[Mux.scala 46:16:@12756.4]
  assign _T_15573 = 6'he == _T_10211_57; // @[Mux.scala 46:19:@12757.4]
  assign _T_15574 = _T_15573 ? _T_9260_13 : _T_15572; // @[Mux.scala 46:16:@12758.4]
  assign _T_15575 = 6'hd == _T_10211_57; // @[Mux.scala 46:19:@12759.4]
  assign _T_15576 = _T_15575 ? _T_9260_12 : _T_15574; // @[Mux.scala 46:16:@12760.4]
  assign _T_15577 = 6'hc == _T_10211_57; // @[Mux.scala 46:19:@12761.4]
  assign _T_15578 = _T_15577 ? _T_9260_11 : _T_15576; // @[Mux.scala 46:16:@12762.4]
  assign _T_15579 = 6'hb == _T_10211_57; // @[Mux.scala 46:19:@12763.4]
  assign _T_15580 = _T_15579 ? _T_9260_10 : _T_15578; // @[Mux.scala 46:16:@12764.4]
  assign _T_15581 = 6'ha == _T_10211_57; // @[Mux.scala 46:19:@12765.4]
  assign _T_15582 = _T_15581 ? _T_9260_9 : _T_15580; // @[Mux.scala 46:16:@12766.4]
  assign _T_15583 = 6'h9 == _T_10211_57; // @[Mux.scala 46:19:@12767.4]
  assign _T_15584 = _T_15583 ? _T_9260_8 : _T_15582; // @[Mux.scala 46:16:@12768.4]
  assign _T_15585 = 6'h8 == _T_10211_57; // @[Mux.scala 46:19:@12769.4]
  assign _T_15586 = _T_15585 ? _T_9260_7 : _T_15584; // @[Mux.scala 46:16:@12770.4]
  assign _T_15587 = 6'h7 == _T_10211_57; // @[Mux.scala 46:19:@12771.4]
  assign _T_15588 = _T_15587 ? _T_9260_6 : _T_15586; // @[Mux.scala 46:16:@12772.4]
  assign _T_15589 = 6'h6 == _T_10211_57; // @[Mux.scala 46:19:@12773.4]
  assign _T_15590 = _T_15589 ? _T_9260_5 : _T_15588; // @[Mux.scala 46:16:@12774.4]
  assign _T_15591 = 6'h5 == _T_10211_57; // @[Mux.scala 46:19:@12775.4]
  assign _T_15592 = _T_15591 ? _T_9260_4 : _T_15590; // @[Mux.scala 46:16:@12776.4]
  assign _T_15593 = 6'h4 == _T_10211_57; // @[Mux.scala 46:19:@12777.4]
  assign _T_15594 = _T_15593 ? _T_9260_3 : _T_15592; // @[Mux.scala 46:16:@12778.4]
  assign _T_15595 = 6'h3 == _T_10211_57; // @[Mux.scala 46:19:@12779.4]
  assign _T_15596 = _T_15595 ? _T_9260_2 : _T_15594; // @[Mux.scala 46:16:@12780.4]
  assign _T_15597 = 6'h2 == _T_10211_57; // @[Mux.scala 46:19:@12781.4]
  assign _T_15598 = _T_15597 ? _T_9260_1 : _T_15596; // @[Mux.scala 46:16:@12782.4]
  assign _T_15599 = 6'h1 == _T_10211_57; // @[Mux.scala 46:19:@12783.4]
  assign _T_15600 = _T_15599 ? _T_9260_0 : _T_15598; // @[Mux.scala 46:16:@12784.4]
  assign _T_15661 = 6'h3b == _T_10211_58; // @[Mux.scala 46:19:@12786.4]
  assign _T_15662 = _T_15661 ? _T_9260_58 : 8'h0; // @[Mux.scala 46:16:@12787.4]
  assign _T_15663 = 6'h3a == _T_10211_58; // @[Mux.scala 46:19:@12788.4]
  assign _T_15664 = _T_15663 ? _T_9260_57 : _T_15662; // @[Mux.scala 46:16:@12789.4]
  assign _T_15665 = 6'h39 == _T_10211_58; // @[Mux.scala 46:19:@12790.4]
  assign _T_15666 = _T_15665 ? _T_9260_56 : _T_15664; // @[Mux.scala 46:16:@12791.4]
  assign _T_15667 = 6'h38 == _T_10211_58; // @[Mux.scala 46:19:@12792.4]
  assign _T_15668 = _T_15667 ? _T_9260_55 : _T_15666; // @[Mux.scala 46:16:@12793.4]
  assign _T_15669 = 6'h37 == _T_10211_58; // @[Mux.scala 46:19:@12794.4]
  assign _T_15670 = _T_15669 ? _T_9260_54 : _T_15668; // @[Mux.scala 46:16:@12795.4]
  assign _T_15671 = 6'h36 == _T_10211_58; // @[Mux.scala 46:19:@12796.4]
  assign _T_15672 = _T_15671 ? _T_9260_53 : _T_15670; // @[Mux.scala 46:16:@12797.4]
  assign _T_15673 = 6'h35 == _T_10211_58; // @[Mux.scala 46:19:@12798.4]
  assign _T_15674 = _T_15673 ? _T_9260_52 : _T_15672; // @[Mux.scala 46:16:@12799.4]
  assign _T_15675 = 6'h34 == _T_10211_58; // @[Mux.scala 46:19:@12800.4]
  assign _T_15676 = _T_15675 ? _T_9260_51 : _T_15674; // @[Mux.scala 46:16:@12801.4]
  assign _T_15677 = 6'h33 == _T_10211_58; // @[Mux.scala 46:19:@12802.4]
  assign _T_15678 = _T_15677 ? _T_9260_50 : _T_15676; // @[Mux.scala 46:16:@12803.4]
  assign _T_15679 = 6'h32 == _T_10211_58; // @[Mux.scala 46:19:@12804.4]
  assign _T_15680 = _T_15679 ? _T_9260_49 : _T_15678; // @[Mux.scala 46:16:@12805.4]
  assign _T_15681 = 6'h31 == _T_10211_58; // @[Mux.scala 46:19:@12806.4]
  assign _T_15682 = _T_15681 ? _T_9260_48 : _T_15680; // @[Mux.scala 46:16:@12807.4]
  assign _T_15683 = 6'h30 == _T_10211_58; // @[Mux.scala 46:19:@12808.4]
  assign _T_15684 = _T_15683 ? _T_9260_47 : _T_15682; // @[Mux.scala 46:16:@12809.4]
  assign _T_15685 = 6'h2f == _T_10211_58; // @[Mux.scala 46:19:@12810.4]
  assign _T_15686 = _T_15685 ? _T_9260_46 : _T_15684; // @[Mux.scala 46:16:@12811.4]
  assign _T_15687 = 6'h2e == _T_10211_58; // @[Mux.scala 46:19:@12812.4]
  assign _T_15688 = _T_15687 ? _T_9260_45 : _T_15686; // @[Mux.scala 46:16:@12813.4]
  assign _T_15689 = 6'h2d == _T_10211_58; // @[Mux.scala 46:19:@12814.4]
  assign _T_15690 = _T_15689 ? _T_9260_44 : _T_15688; // @[Mux.scala 46:16:@12815.4]
  assign _T_15691 = 6'h2c == _T_10211_58; // @[Mux.scala 46:19:@12816.4]
  assign _T_15692 = _T_15691 ? _T_9260_43 : _T_15690; // @[Mux.scala 46:16:@12817.4]
  assign _T_15693 = 6'h2b == _T_10211_58; // @[Mux.scala 46:19:@12818.4]
  assign _T_15694 = _T_15693 ? _T_9260_42 : _T_15692; // @[Mux.scala 46:16:@12819.4]
  assign _T_15695 = 6'h2a == _T_10211_58; // @[Mux.scala 46:19:@12820.4]
  assign _T_15696 = _T_15695 ? _T_9260_41 : _T_15694; // @[Mux.scala 46:16:@12821.4]
  assign _T_15697 = 6'h29 == _T_10211_58; // @[Mux.scala 46:19:@12822.4]
  assign _T_15698 = _T_15697 ? _T_9260_40 : _T_15696; // @[Mux.scala 46:16:@12823.4]
  assign _T_15699 = 6'h28 == _T_10211_58; // @[Mux.scala 46:19:@12824.4]
  assign _T_15700 = _T_15699 ? _T_9260_39 : _T_15698; // @[Mux.scala 46:16:@12825.4]
  assign _T_15701 = 6'h27 == _T_10211_58; // @[Mux.scala 46:19:@12826.4]
  assign _T_15702 = _T_15701 ? _T_9260_38 : _T_15700; // @[Mux.scala 46:16:@12827.4]
  assign _T_15703 = 6'h26 == _T_10211_58; // @[Mux.scala 46:19:@12828.4]
  assign _T_15704 = _T_15703 ? _T_9260_37 : _T_15702; // @[Mux.scala 46:16:@12829.4]
  assign _T_15705 = 6'h25 == _T_10211_58; // @[Mux.scala 46:19:@12830.4]
  assign _T_15706 = _T_15705 ? _T_9260_36 : _T_15704; // @[Mux.scala 46:16:@12831.4]
  assign _T_15707 = 6'h24 == _T_10211_58; // @[Mux.scala 46:19:@12832.4]
  assign _T_15708 = _T_15707 ? _T_9260_35 : _T_15706; // @[Mux.scala 46:16:@12833.4]
  assign _T_15709 = 6'h23 == _T_10211_58; // @[Mux.scala 46:19:@12834.4]
  assign _T_15710 = _T_15709 ? _T_9260_34 : _T_15708; // @[Mux.scala 46:16:@12835.4]
  assign _T_15711 = 6'h22 == _T_10211_58; // @[Mux.scala 46:19:@12836.4]
  assign _T_15712 = _T_15711 ? _T_9260_33 : _T_15710; // @[Mux.scala 46:16:@12837.4]
  assign _T_15713 = 6'h21 == _T_10211_58; // @[Mux.scala 46:19:@12838.4]
  assign _T_15714 = _T_15713 ? _T_9260_32 : _T_15712; // @[Mux.scala 46:16:@12839.4]
  assign _T_15715 = 6'h20 == _T_10211_58; // @[Mux.scala 46:19:@12840.4]
  assign _T_15716 = _T_15715 ? _T_9260_31 : _T_15714; // @[Mux.scala 46:16:@12841.4]
  assign _T_15717 = 6'h1f == _T_10211_58; // @[Mux.scala 46:19:@12842.4]
  assign _T_15718 = _T_15717 ? _T_9260_30 : _T_15716; // @[Mux.scala 46:16:@12843.4]
  assign _T_15719 = 6'h1e == _T_10211_58; // @[Mux.scala 46:19:@12844.4]
  assign _T_15720 = _T_15719 ? _T_9260_29 : _T_15718; // @[Mux.scala 46:16:@12845.4]
  assign _T_15721 = 6'h1d == _T_10211_58; // @[Mux.scala 46:19:@12846.4]
  assign _T_15722 = _T_15721 ? _T_9260_28 : _T_15720; // @[Mux.scala 46:16:@12847.4]
  assign _T_15723 = 6'h1c == _T_10211_58; // @[Mux.scala 46:19:@12848.4]
  assign _T_15724 = _T_15723 ? _T_9260_27 : _T_15722; // @[Mux.scala 46:16:@12849.4]
  assign _T_15725 = 6'h1b == _T_10211_58; // @[Mux.scala 46:19:@12850.4]
  assign _T_15726 = _T_15725 ? _T_9260_26 : _T_15724; // @[Mux.scala 46:16:@12851.4]
  assign _T_15727 = 6'h1a == _T_10211_58; // @[Mux.scala 46:19:@12852.4]
  assign _T_15728 = _T_15727 ? _T_9260_25 : _T_15726; // @[Mux.scala 46:16:@12853.4]
  assign _T_15729 = 6'h19 == _T_10211_58; // @[Mux.scala 46:19:@12854.4]
  assign _T_15730 = _T_15729 ? _T_9260_24 : _T_15728; // @[Mux.scala 46:16:@12855.4]
  assign _T_15731 = 6'h18 == _T_10211_58; // @[Mux.scala 46:19:@12856.4]
  assign _T_15732 = _T_15731 ? _T_9260_23 : _T_15730; // @[Mux.scala 46:16:@12857.4]
  assign _T_15733 = 6'h17 == _T_10211_58; // @[Mux.scala 46:19:@12858.4]
  assign _T_15734 = _T_15733 ? _T_9260_22 : _T_15732; // @[Mux.scala 46:16:@12859.4]
  assign _T_15735 = 6'h16 == _T_10211_58; // @[Mux.scala 46:19:@12860.4]
  assign _T_15736 = _T_15735 ? _T_9260_21 : _T_15734; // @[Mux.scala 46:16:@12861.4]
  assign _T_15737 = 6'h15 == _T_10211_58; // @[Mux.scala 46:19:@12862.4]
  assign _T_15738 = _T_15737 ? _T_9260_20 : _T_15736; // @[Mux.scala 46:16:@12863.4]
  assign _T_15739 = 6'h14 == _T_10211_58; // @[Mux.scala 46:19:@12864.4]
  assign _T_15740 = _T_15739 ? _T_9260_19 : _T_15738; // @[Mux.scala 46:16:@12865.4]
  assign _T_15741 = 6'h13 == _T_10211_58; // @[Mux.scala 46:19:@12866.4]
  assign _T_15742 = _T_15741 ? _T_9260_18 : _T_15740; // @[Mux.scala 46:16:@12867.4]
  assign _T_15743 = 6'h12 == _T_10211_58; // @[Mux.scala 46:19:@12868.4]
  assign _T_15744 = _T_15743 ? _T_9260_17 : _T_15742; // @[Mux.scala 46:16:@12869.4]
  assign _T_15745 = 6'h11 == _T_10211_58; // @[Mux.scala 46:19:@12870.4]
  assign _T_15746 = _T_15745 ? _T_9260_16 : _T_15744; // @[Mux.scala 46:16:@12871.4]
  assign _T_15747 = 6'h10 == _T_10211_58; // @[Mux.scala 46:19:@12872.4]
  assign _T_15748 = _T_15747 ? _T_9260_15 : _T_15746; // @[Mux.scala 46:16:@12873.4]
  assign _T_15749 = 6'hf == _T_10211_58; // @[Mux.scala 46:19:@12874.4]
  assign _T_15750 = _T_15749 ? _T_9260_14 : _T_15748; // @[Mux.scala 46:16:@12875.4]
  assign _T_15751 = 6'he == _T_10211_58; // @[Mux.scala 46:19:@12876.4]
  assign _T_15752 = _T_15751 ? _T_9260_13 : _T_15750; // @[Mux.scala 46:16:@12877.4]
  assign _T_15753 = 6'hd == _T_10211_58; // @[Mux.scala 46:19:@12878.4]
  assign _T_15754 = _T_15753 ? _T_9260_12 : _T_15752; // @[Mux.scala 46:16:@12879.4]
  assign _T_15755 = 6'hc == _T_10211_58; // @[Mux.scala 46:19:@12880.4]
  assign _T_15756 = _T_15755 ? _T_9260_11 : _T_15754; // @[Mux.scala 46:16:@12881.4]
  assign _T_15757 = 6'hb == _T_10211_58; // @[Mux.scala 46:19:@12882.4]
  assign _T_15758 = _T_15757 ? _T_9260_10 : _T_15756; // @[Mux.scala 46:16:@12883.4]
  assign _T_15759 = 6'ha == _T_10211_58; // @[Mux.scala 46:19:@12884.4]
  assign _T_15760 = _T_15759 ? _T_9260_9 : _T_15758; // @[Mux.scala 46:16:@12885.4]
  assign _T_15761 = 6'h9 == _T_10211_58; // @[Mux.scala 46:19:@12886.4]
  assign _T_15762 = _T_15761 ? _T_9260_8 : _T_15760; // @[Mux.scala 46:16:@12887.4]
  assign _T_15763 = 6'h8 == _T_10211_58; // @[Mux.scala 46:19:@12888.4]
  assign _T_15764 = _T_15763 ? _T_9260_7 : _T_15762; // @[Mux.scala 46:16:@12889.4]
  assign _T_15765 = 6'h7 == _T_10211_58; // @[Mux.scala 46:19:@12890.4]
  assign _T_15766 = _T_15765 ? _T_9260_6 : _T_15764; // @[Mux.scala 46:16:@12891.4]
  assign _T_15767 = 6'h6 == _T_10211_58; // @[Mux.scala 46:19:@12892.4]
  assign _T_15768 = _T_15767 ? _T_9260_5 : _T_15766; // @[Mux.scala 46:16:@12893.4]
  assign _T_15769 = 6'h5 == _T_10211_58; // @[Mux.scala 46:19:@12894.4]
  assign _T_15770 = _T_15769 ? _T_9260_4 : _T_15768; // @[Mux.scala 46:16:@12895.4]
  assign _T_15771 = 6'h4 == _T_10211_58; // @[Mux.scala 46:19:@12896.4]
  assign _T_15772 = _T_15771 ? _T_9260_3 : _T_15770; // @[Mux.scala 46:16:@12897.4]
  assign _T_15773 = 6'h3 == _T_10211_58; // @[Mux.scala 46:19:@12898.4]
  assign _T_15774 = _T_15773 ? _T_9260_2 : _T_15772; // @[Mux.scala 46:16:@12899.4]
  assign _T_15775 = 6'h2 == _T_10211_58; // @[Mux.scala 46:19:@12900.4]
  assign _T_15776 = _T_15775 ? _T_9260_1 : _T_15774; // @[Mux.scala 46:16:@12901.4]
  assign _T_15777 = 6'h1 == _T_10211_58; // @[Mux.scala 46:19:@12902.4]
  assign _T_15778 = _T_15777 ? _T_9260_0 : _T_15776; // @[Mux.scala 46:16:@12903.4]
  assign _T_15840 = 6'h3c == _T_10211_59; // @[Mux.scala 46:19:@12905.4]
  assign _T_15841 = _T_15840 ? _T_9260_59 : 8'h0; // @[Mux.scala 46:16:@12906.4]
  assign _T_15842 = 6'h3b == _T_10211_59; // @[Mux.scala 46:19:@12907.4]
  assign _T_15843 = _T_15842 ? _T_9260_58 : _T_15841; // @[Mux.scala 46:16:@12908.4]
  assign _T_15844 = 6'h3a == _T_10211_59; // @[Mux.scala 46:19:@12909.4]
  assign _T_15845 = _T_15844 ? _T_9260_57 : _T_15843; // @[Mux.scala 46:16:@12910.4]
  assign _T_15846 = 6'h39 == _T_10211_59; // @[Mux.scala 46:19:@12911.4]
  assign _T_15847 = _T_15846 ? _T_9260_56 : _T_15845; // @[Mux.scala 46:16:@12912.4]
  assign _T_15848 = 6'h38 == _T_10211_59; // @[Mux.scala 46:19:@12913.4]
  assign _T_15849 = _T_15848 ? _T_9260_55 : _T_15847; // @[Mux.scala 46:16:@12914.4]
  assign _T_15850 = 6'h37 == _T_10211_59; // @[Mux.scala 46:19:@12915.4]
  assign _T_15851 = _T_15850 ? _T_9260_54 : _T_15849; // @[Mux.scala 46:16:@12916.4]
  assign _T_15852 = 6'h36 == _T_10211_59; // @[Mux.scala 46:19:@12917.4]
  assign _T_15853 = _T_15852 ? _T_9260_53 : _T_15851; // @[Mux.scala 46:16:@12918.4]
  assign _T_15854 = 6'h35 == _T_10211_59; // @[Mux.scala 46:19:@12919.4]
  assign _T_15855 = _T_15854 ? _T_9260_52 : _T_15853; // @[Mux.scala 46:16:@12920.4]
  assign _T_15856 = 6'h34 == _T_10211_59; // @[Mux.scala 46:19:@12921.4]
  assign _T_15857 = _T_15856 ? _T_9260_51 : _T_15855; // @[Mux.scala 46:16:@12922.4]
  assign _T_15858 = 6'h33 == _T_10211_59; // @[Mux.scala 46:19:@12923.4]
  assign _T_15859 = _T_15858 ? _T_9260_50 : _T_15857; // @[Mux.scala 46:16:@12924.4]
  assign _T_15860 = 6'h32 == _T_10211_59; // @[Mux.scala 46:19:@12925.4]
  assign _T_15861 = _T_15860 ? _T_9260_49 : _T_15859; // @[Mux.scala 46:16:@12926.4]
  assign _T_15862 = 6'h31 == _T_10211_59; // @[Mux.scala 46:19:@12927.4]
  assign _T_15863 = _T_15862 ? _T_9260_48 : _T_15861; // @[Mux.scala 46:16:@12928.4]
  assign _T_15864 = 6'h30 == _T_10211_59; // @[Mux.scala 46:19:@12929.4]
  assign _T_15865 = _T_15864 ? _T_9260_47 : _T_15863; // @[Mux.scala 46:16:@12930.4]
  assign _T_15866 = 6'h2f == _T_10211_59; // @[Mux.scala 46:19:@12931.4]
  assign _T_15867 = _T_15866 ? _T_9260_46 : _T_15865; // @[Mux.scala 46:16:@12932.4]
  assign _T_15868 = 6'h2e == _T_10211_59; // @[Mux.scala 46:19:@12933.4]
  assign _T_15869 = _T_15868 ? _T_9260_45 : _T_15867; // @[Mux.scala 46:16:@12934.4]
  assign _T_15870 = 6'h2d == _T_10211_59; // @[Mux.scala 46:19:@12935.4]
  assign _T_15871 = _T_15870 ? _T_9260_44 : _T_15869; // @[Mux.scala 46:16:@12936.4]
  assign _T_15872 = 6'h2c == _T_10211_59; // @[Mux.scala 46:19:@12937.4]
  assign _T_15873 = _T_15872 ? _T_9260_43 : _T_15871; // @[Mux.scala 46:16:@12938.4]
  assign _T_15874 = 6'h2b == _T_10211_59; // @[Mux.scala 46:19:@12939.4]
  assign _T_15875 = _T_15874 ? _T_9260_42 : _T_15873; // @[Mux.scala 46:16:@12940.4]
  assign _T_15876 = 6'h2a == _T_10211_59; // @[Mux.scala 46:19:@12941.4]
  assign _T_15877 = _T_15876 ? _T_9260_41 : _T_15875; // @[Mux.scala 46:16:@12942.4]
  assign _T_15878 = 6'h29 == _T_10211_59; // @[Mux.scala 46:19:@12943.4]
  assign _T_15879 = _T_15878 ? _T_9260_40 : _T_15877; // @[Mux.scala 46:16:@12944.4]
  assign _T_15880 = 6'h28 == _T_10211_59; // @[Mux.scala 46:19:@12945.4]
  assign _T_15881 = _T_15880 ? _T_9260_39 : _T_15879; // @[Mux.scala 46:16:@12946.4]
  assign _T_15882 = 6'h27 == _T_10211_59; // @[Mux.scala 46:19:@12947.4]
  assign _T_15883 = _T_15882 ? _T_9260_38 : _T_15881; // @[Mux.scala 46:16:@12948.4]
  assign _T_15884 = 6'h26 == _T_10211_59; // @[Mux.scala 46:19:@12949.4]
  assign _T_15885 = _T_15884 ? _T_9260_37 : _T_15883; // @[Mux.scala 46:16:@12950.4]
  assign _T_15886 = 6'h25 == _T_10211_59; // @[Mux.scala 46:19:@12951.4]
  assign _T_15887 = _T_15886 ? _T_9260_36 : _T_15885; // @[Mux.scala 46:16:@12952.4]
  assign _T_15888 = 6'h24 == _T_10211_59; // @[Mux.scala 46:19:@12953.4]
  assign _T_15889 = _T_15888 ? _T_9260_35 : _T_15887; // @[Mux.scala 46:16:@12954.4]
  assign _T_15890 = 6'h23 == _T_10211_59; // @[Mux.scala 46:19:@12955.4]
  assign _T_15891 = _T_15890 ? _T_9260_34 : _T_15889; // @[Mux.scala 46:16:@12956.4]
  assign _T_15892 = 6'h22 == _T_10211_59; // @[Mux.scala 46:19:@12957.4]
  assign _T_15893 = _T_15892 ? _T_9260_33 : _T_15891; // @[Mux.scala 46:16:@12958.4]
  assign _T_15894 = 6'h21 == _T_10211_59; // @[Mux.scala 46:19:@12959.4]
  assign _T_15895 = _T_15894 ? _T_9260_32 : _T_15893; // @[Mux.scala 46:16:@12960.4]
  assign _T_15896 = 6'h20 == _T_10211_59; // @[Mux.scala 46:19:@12961.4]
  assign _T_15897 = _T_15896 ? _T_9260_31 : _T_15895; // @[Mux.scala 46:16:@12962.4]
  assign _T_15898 = 6'h1f == _T_10211_59; // @[Mux.scala 46:19:@12963.4]
  assign _T_15899 = _T_15898 ? _T_9260_30 : _T_15897; // @[Mux.scala 46:16:@12964.4]
  assign _T_15900 = 6'h1e == _T_10211_59; // @[Mux.scala 46:19:@12965.4]
  assign _T_15901 = _T_15900 ? _T_9260_29 : _T_15899; // @[Mux.scala 46:16:@12966.4]
  assign _T_15902 = 6'h1d == _T_10211_59; // @[Mux.scala 46:19:@12967.4]
  assign _T_15903 = _T_15902 ? _T_9260_28 : _T_15901; // @[Mux.scala 46:16:@12968.4]
  assign _T_15904 = 6'h1c == _T_10211_59; // @[Mux.scala 46:19:@12969.4]
  assign _T_15905 = _T_15904 ? _T_9260_27 : _T_15903; // @[Mux.scala 46:16:@12970.4]
  assign _T_15906 = 6'h1b == _T_10211_59; // @[Mux.scala 46:19:@12971.4]
  assign _T_15907 = _T_15906 ? _T_9260_26 : _T_15905; // @[Mux.scala 46:16:@12972.4]
  assign _T_15908 = 6'h1a == _T_10211_59; // @[Mux.scala 46:19:@12973.4]
  assign _T_15909 = _T_15908 ? _T_9260_25 : _T_15907; // @[Mux.scala 46:16:@12974.4]
  assign _T_15910 = 6'h19 == _T_10211_59; // @[Mux.scala 46:19:@12975.4]
  assign _T_15911 = _T_15910 ? _T_9260_24 : _T_15909; // @[Mux.scala 46:16:@12976.4]
  assign _T_15912 = 6'h18 == _T_10211_59; // @[Mux.scala 46:19:@12977.4]
  assign _T_15913 = _T_15912 ? _T_9260_23 : _T_15911; // @[Mux.scala 46:16:@12978.4]
  assign _T_15914 = 6'h17 == _T_10211_59; // @[Mux.scala 46:19:@12979.4]
  assign _T_15915 = _T_15914 ? _T_9260_22 : _T_15913; // @[Mux.scala 46:16:@12980.4]
  assign _T_15916 = 6'h16 == _T_10211_59; // @[Mux.scala 46:19:@12981.4]
  assign _T_15917 = _T_15916 ? _T_9260_21 : _T_15915; // @[Mux.scala 46:16:@12982.4]
  assign _T_15918 = 6'h15 == _T_10211_59; // @[Mux.scala 46:19:@12983.4]
  assign _T_15919 = _T_15918 ? _T_9260_20 : _T_15917; // @[Mux.scala 46:16:@12984.4]
  assign _T_15920 = 6'h14 == _T_10211_59; // @[Mux.scala 46:19:@12985.4]
  assign _T_15921 = _T_15920 ? _T_9260_19 : _T_15919; // @[Mux.scala 46:16:@12986.4]
  assign _T_15922 = 6'h13 == _T_10211_59; // @[Mux.scala 46:19:@12987.4]
  assign _T_15923 = _T_15922 ? _T_9260_18 : _T_15921; // @[Mux.scala 46:16:@12988.4]
  assign _T_15924 = 6'h12 == _T_10211_59; // @[Mux.scala 46:19:@12989.4]
  assign _T_15925 = _T_15924 ? _T_9260_17 : _T_15923; // @[Mux.scala 46:16:@12990.4]
  assign _T_15926 = 6'h11 == _T_10211_59; // @[Mux.scala 46:19:@12991.4]
  assign _T_15927 = _T_15926 ? _T_9260_16 : _T_15925; // @[Mux.scala 46:16:@12992.4]
  assign _T_15928 = 6'h10 == _T_10211_59; // @[Mux.scala 46:19:@12993.4]
  assign _T_15929 = _T_15928 ? _T_9260_15 : _T_15927; // @[Mux.scala 46:16:@12994.4]
  assign _T_15930 = 6'hf == _T_10211_59; // @[Mux.scala 46:19:@12995.4]
  assign _T_15931 = _T_15930 ? _T_9260_14 : _T_15929; // @[Mux.scala 46:16:@12996.4]
  assign _T_15932 = 6'he == _T_10211_59; // @[Mux.scala 46:19:@12997.4]
  assign _T_15933 = _T_15932 ? _T_9260_13 : _T_15931; // @[Mux.scala 46:16:@12998.4]
  assign _T_15934 = 6'hd == _T_10211_59; // @[Mux.scala 46:19:@12999.4]
  assign _T_15935 = _T_15934 ? _T_9260_12 : _T_15933; // @[Mux.scala 46:16:@13000.4]
  assign _T_15936 = 6'hc == _T_10211_59; // @[Mux.scala 46:19:@13001.4]
  assign _T_15937 = _T_15936 ? _T_9260_11 : _T_15935; // @[Mux.scala 46:16:@13002.4]
  assign _T_15938 = 6'hb == _T_10211_59; // @[Mux.scala 46:19:@13003.4]
  assign _T_15939 = _T_15938 ? _T_9260_10 : _T_15937; // @[Mux.scala 46:16:@13004.4]
  assign _T_15940 = 6'ha == _T_10211_59; // @[Mux.scala 46:19:@13005.4]
  assign _T_15941 = _T_15940 ? _T_9260_9 : _T_15939; // @[Mux.scala 46:16:@13006.4]
  assign _T_15942 = 6'h9 == _T_10211_59; // @[Mux.scala 46:19:@13007.4]
  assign _T_15943 = _T_15942 ? _T_9260_8 : _T_15941; // @[Mux.scala 46:16:@13008.4]
  assign _T_15944 = 6'h8 == _T_10211_59; // @[Mux.scala 46:19:@13009.4]
  assign _T_15945 = _T_15944 ? _T_9260_7 : _T_15943; // @[Mux.scala 46:16:@13010.4]
  assign _T_15946 = 6'h7 == _T_10211_59; // @[Mux.scala 46:19:@13011.4]
  assign _T_15947 = _T_15946 ? _T_9260_6 : _T_15945; // @[Mux.scala 46:16:@13012.4]
  assign _T_15948 = 6'h6 == _T_10211_59; // @[Mux.scala 46:19:@13013.4]
  assign _T_15949 = _T_15948 ? _T_9260_5 : _T_15947; // @[Mux.scala 46:16:@13014.4]
  assign _T_15950 = 6'h5 == _T_10211_59; // @[Mux.scala 46:19:@13015.4]
  assign _T_15951 = _T_15950 ? _T_9260_4 : _T_15949; // @[Mux.scala 46:16:@13016.4]
  assign _T_15952 = 6'h4 == _T_10211_59; // @[Mux.scala 46:19:@13017.4]
  assign _T_15953 = _T_15952 ? _T_9260_3 : _T_15951; // @[Mux.scala 46:16:@13018.4]
  assign _T_15954 = 6'h3 == _T_10211_59; // @[Mux.scala 46:19:@13019.4]
  assign _T_15955 = _T_15954 ? _T_9260_2 : _T_15953; // @[Mux.scala 46:16:@13020.4]
  assign _T_15956 = 6'h2 == _T_10211_59; // @[Mux.scala 46:19:@13021.4]
  assign _T_15957 = _T_15956 ? _T_9260_1 : _T_15955; // @[Mux.scala 46:16:@13022.4]
  assign _T_15958 = 6'h1 == _T_10211_59; // @[Mux.scala 46:19:@13023.4]
  assign _T_15959 = _T_15958 ? _T_9260_0 : _T_15957; // @[Mux.scala 46:16:@13024.4]
  assign _T_16022 = 6'h3d == _T_10211_60; // @[Mux.scala 46:19:@13026.4]
  assign _T_16023 = _T_16022 ? _T_9260_60 : 8'h0; // @[Mux.scala 46:16:@13027.4]
  assign _T_16024 = 6'h3c == _T_10211_60; // @[Mux.scala 46:19:@13028.4]
  assign _T_16025 = _T_16024 ? _T_9260_59 : _T_16023; // @[Mux.scala 46:16:@13029.4]
  assign _T_16026 = 6'h3b == _T_10211_60; // @[Mux.scala 46:19:@13030.4]
  assign _T_16027 = _T_16026 ? _T_9260_58 : _T_16025; // @[Mux.scala 46:16:@13031.4]
  assign _T_16028 = 6'h3a == _T_10211_60; // @[Mux.scala 46:19:@13032.4]
  assign _T_16029 = _T_16028 ? _T_9260_57 : _T_16027; // @[Mux.scala 46:16:@13033.4]
  assign _T_16030 = 6'h39 == _T_10211_60; // @[Mux.scala 46:19:@13034.4]
  assign _T_16031 = _T_16030 ? _T_9260_56 : _T_16029; // @[Mux.scala 46:16:@13035.4]
  assign _T_16032 = 6'h38 == _T_10211_60; // @[Mux.scala 46:19:@13036.4]
  assign _T_16033 = _T_16032 ? _T_9260_55 : _T_16031; // @[Mux.scala 46:16:@13037.4]
  assign _T_16034 = 6'h37 == _T_10211_60; // @[Mux.scala 46:19:@13038.4]
  assign _T_16035 = _T_16034 ? _T_9260_54 : _T_16033; // @[Mux.scala 46:16:@13039.4]
  assign _T_16036 = 6'h36 == _T_10211_60; // @[Mux.scala 46:19:@13040.4]
  assign _T_16037 = _T_16036 ? _T_9260_53 : _T_16035; // @[Mux.scala 46:16:@13041.4]
  assign _T_16038 = 6'h35 == _T_10211_60; // @[Mux.scala 46:19:@13042.4]
  assign _T_16039 = _T_16038 ? _T_9260_52 : _T_16037; // @[Mux.scala 46:16:@13043.4]
  assign _T_16040 = 6'h34 == _T_10211_60; // @[Mux.scala 46:19:@13044.4]
  assign _T_16041 = _T_16040 ? _T_9260_51 : _T_16039; // @[Mux.scala 46:16:@13045.4]
  assign _T_16042 = 6'h33 == _T_10211_60; // @[Mux.scala 46:19:@13046.4]
  assign _T_16043 = _T_16042 ? _T_9260_50 : _T_16041; // @[Mux.scala 46:16:@13047.4]
  assign _T_16044 = 6'h32 == _T_10211_60; // @[Mux.scala 46:19:@13048.4]
  assign _T_16045 = _T_16044 ? _T_9260_49 : _T_16043; // @[Mux.scala 46:16:@13049.4]
  assign _T_16046 = 6'h31 == _T_10211_60; // @[Mux.scala 46:19:@13050.4]
  assign _T_16047 = _T_16046 ? _T_9260_48 : _T_16045; // @[Mux.scala 46:16:@13051.4]
  assign _T_16048 = 6'h30 == _T_10211_60; // @[Mux.scala 46:19:@13052.4]
  assign _T_16049 = _T_16048 ? _T_9260_47 : _T_16047; // @[Mux.scala 46:16:@13053.4]
  assign _T_16050 = 6'h2f == _T_10211_60; // @[Mux.scala 46:19:@13054.4]
  assign _T_16051 = _T_16050 ? _T_9260_46 : _T_16049; // @[Mux.scala 46:16:@13055.4]
  assign _T_16052 = 6'h2e == _T_10211_60; // @[Mux.scala 46:19:@13056.4]
  assign _T_16053 = _T_16052 ? _T_9260_45 : _T_16051; // @[Mux.scala 46:16:@13057.4]
  assign _T_16054 = 6'h2d == _T_10211_60; // @[Mux.scala 46:19:@13058.4]
  assign _T_16055 = _T_16054 ? _T_9260_44 : _T_16053; // @[Mux.scala 46:16:@13059.4]
  assign _T_16056 = 6'h2c == _T_10211_60; // @[Mux.scala 46:19:@13060.4]
  assign _T_16057 = _T_16056 ? _T_9260_43 : _T_16055; // @[Mux.scala 46:16:@13061.4]
  assign _T_16058 = 6'h2b == _T_10211_60; // @[Mux.scala 46:19:@13062.4]
  assign _T_16059 = _T_16058 ? _T_9260_42 : _T_16057; // @[Mux.scala 46:16:@13063.4]
  assign _T_16060 = 6'h2a == _T_10211_60; // @[Mux.scala 46:19:@13064.4]
  assign _T_16061 = _T_16060 ? _T_9260_41 : _T_16059; // @[Mux.scala 46:16:@13065.4]
  assign _T_16062 = 6'h29 == _T_10211_60; // @[Mux.scala 46:19:@13066.4]
  assign _T_16063 = _T_16062 ? _T_9260_40 : _T_16061; // @[Mux.scala 46:16:@13067.4]
  assign _T_16064 = 6'h28 == _T_10211_60; // @[Mux.scala 46:19:@13068.4]
  assign _T_16065 = _T_16064 ? _T_9260_39 : _T_16063; // @[Mux.scala 46:16:@13069.4]
  assign _T_16066 = 6'h27 == _T_10211_60; // @[Mux.scala 46:19:@13070.4]
  assign _T_16067 = _T_16066 ? _T_9260_38 : _T_16065; // @[Mux.scala 46:16:@13071.4]
  assign _T_16068 = 6'h26 == _T_10211_60; // @[Mux.scala 46:19:@13072.4]
  assign _T_16069 = _T_16068 ? _T_9260_37 : _T_16067; // @[Mux.scala 46:16:@13073.4]
  assign _T_16070 = 6'h25 == _T_10211_60; // @[Mux.scala 46:19:@13074.4]
  assign _T_16071 = _T_16070 ? _T_9260_36 : _T_16069; // @[Mux.scala 46:16:@13075.4]
  assign _T_16072 = 6'h24 == _T_10211_60; // @[Mux.scala 46:19:@13076.4]
  assign _T_16073 = _T_16072 ? _T_9260_35 : _T_16071; // @[Mux.scala 46:16:@13077.4]
  assign _T_16074 = 6'h23 == _T_10211_60; // @[Mux.scala 46:19:@13078.4]
  assign _T_16075 = _T_16074 ? _T_9260_34 : _T_16073; // @[Mux.scala 46:16:@13079.4]
  assign _T_16076 = 6'h22 == _T_10211_60; // @[Mux.scala 46:19:@13080.4]
  assign _T_16077 = _T_16076 ? _T_9260_33 : _T_16075; // @[Mux.scala 46:16:@13081.4]
  assign _T_16078 = 6'h21 == _T_10211_60; // @[Mux.scala 46:19:@13082.4]
  assign _T_16079 = _T_16078 ? _T_9260_32 : _T_16077; // @[Mux.scala 46:16:@13083.4]
  assign _T_16080 = 6'h20 == _T_10211_60; // @[Mux.scala 46:19:@13084.4]
  assign _T_16081 = _T_16080 ? _T_9260_31 : _T_16079; // @[Mux.scala 46:16:@13085.4]
  assign _T_16082 = 6'h1f == _T_10211_60; // @[Mux.scala 46:19:@13086.4]
  assign _T_16083 = _T_16082 ? _T_9260_30 : _T_16081; // @[Mux.scala 46:16:@13087.4]
  assign _T_16084 = 6'h1e == _T_10211_60; // @[Mux.scala 46:19:@13088.4]
  assign _T_16085 = _T_16084 ? _T_9260_29 : _T_16083; // @[Mux.scala 46:16:@13089.4]
  assign _T_16086 = 6'h1d == _T_10211_60; // @[Mux.scala 46:19:@13090.4]
  assign _T_16087 = _T_16086 ? _T_9260_28 : _T_16085; // @[Mux.scala 46:16:@13091.4]
  assign _T_16088 = 6'h1c == _T_10211_60; // @[Mux.scala 46:19:@13092.4]
  assign _T_16089 = _T_16088 ? _T_9260_27 : _T_16087; // @[Mux.scala 46:16:@13093.4]
  assign _T_16090 = 6'h1b == _T_10211_60; // @[Mux.scala 46:19:@13094.4]
  assign _T_16091 = _T_16090 ? _T_9260_26 : _T_16089; // @[Mux.scala 46:16:@13095.4]
  assign _T_16092 = 6'h1a == _T_10211_60; // @[Mux.scala 46:19:@13096.4]
  assign _T_16093 = _T_16092 ? _T_9260_25 : _T_16091; // @[Mux.scala 46:16:@13097.4]
  assign _T_16094 = 6'h19 == _T_10211_60; // @[Mux.scala 46:19:@13098.4]
  assign _T_16095 = _T_16094 ? _T_9260_24 : _T_16093; // @[Mux.scala 46:16:@13099.4]
  assign _T_16096 = 6'h18 == _T_10211_60; // @[Mux.scala 46:19:@13100.4]
  assign _T_16097 = _T_16096 ? _T_9260_23 : _T_16095; // @[Mux.scala 46:16:@13101.4]
  assign _T_16098 = 6'h17 == _T_10211_60; // @[Mux.scala 46:19:@13102.4]
  assign _T_16099 = _T_16098 ? _T_9260_22 : _T_16097; // @[Mux.scala 46:16:@13103.4]
  assign _T_16100 = 6'h16 == _T_10211_60; // @[Mux.scala 46:19:@13104.4]
  assign _T_16101 = _T_16100 ? _T_9260_21 : _T_16099; // @[Mux.scala 46:16:@13105.4]
  assign _T_16102 = 6'h15 == _T_10211_60; // @[Mux.scala 46:19:@13106.4]
  assign _T_16103 = _T_16102 ? _T_9260_20 : _T_16101; // @[Mux.scala 46:16:@13107.4]
  assign _T_16104 = 6'h14 == _T_10211_60; // @[Mux.scala 46:19:@13108.4]
  assign _T_16105 = _T_16104 ? _T_9260_19 : _T_16103; // @[Mux.scala 46:16:@13109.4]
  assign _T_16106 = 6'h13 == _T_10211_60; // @[Mux.scala 46:19:@13110.4]
  assign _T_16107 = _T_16106 ? _T_9260_18 : _T_16105; // @[Mux.scala 46:16:@13111.4]
  assign _T_16108 = 6'h12 == _T_10211_60; // @[Mux.scala 46:19:@13112.4]
  assign _T_16109 = _T_16108 ? _T_9260_17 : _T_16107; // @[Mux.scala 46:16:@13113.4]
  assign _T_16110 = 6'h11 == _T_10211_60; // @[Mux.scala 46:19:@13114.4]
  assign _T_16111 = _T_16110 ? _T_9260_16 : _T_16109; // @[Mux.scala 46:16:@13115.4]
  assign _T_16112 = 6'h10 == _T_10211_60; // @[Mux.scala 46:19:@13116.4]
  assign _T_16113 = _T_16112 ? _T_9260_15 : _T_16111; // @[Mux.scala 46:16:@13117.4]
  assign _T_16114 = 6'hf == _T_10211_60; // @[Mux.scala 46:19:@13118.4]
  assign _T_16115 = _T_16114 ? _T_9260_14 : _T_16113; // @[Mux.scala 46:16:@13119.4]
  assign _T_16116 = 6'he == _T_10211_60; // @[Mux.scala 46:19:@13120.4]
  assign _T_16117 = _T_16116 ? _T_9260_13 : _T_16115; // @[Mux.scala 46:16:@13121.4]
  assign _T_16118 = 6'hd == _T_10211_60; // @[Mux.scala 46:19:@13122.4]
  assign _T_16119 = _T_16118 ? _T_9260_12 : _T_16117; // @[Mux.scala 46:16:@13123.4]
  assign _T_16120 = 6'hc == _T_10211_60; // @[Mux.scala 46:19:@13124.4]
  assign _T_16121 = _T_16120 ? _T_9260_11 : _T_16119; // @[Mux.scala 46:16:@13125.4]
  assign _T_16122 = 6'hb == _T_10211_60; // @[Mux.scala 46:19:@13126.4]
  assign _T_16123 = _T_16122 ? _T_9260_10 : _T_16121; // @[Mux.scala 46:16:@13127.4]
  assign _T_16124 = 6'ha == _T_10211_60; // @[Mux.scala 46:19:@13128.4]
  assign _T_16125 = _T_16124 ? _T_9260_9 : _T_16123; // @[Mux.scala 46:16:@13129.4]
  assign _T_16126 = 6'h9 == _T_10211_60; // @[Mux.scala 46:19:@13130.4]
  assign _T_16127 = _T_16126 ? _T_9260_8 : _T_16125; // @[Mux.scala 46:16:@13131.4]
  assign _T_16128 = 6'h8 == _T_10211_60; // @[Mux.scala 46:19:@13132.4]
  assign _T_16129 = _T_16128 ? _T_9260_7 : _T_16127; // @[Mux.scala 46:16:@13133.4]
  assign _T_16130 = 6'h7 == _T_10211_60; // @[Mux.scala 46:19:@13134.4]
  assign _T_16131 = _T_16130 ? _T_9260_6 : _T_16129; // @[Mux.scala 46:16:@13135.4]
  assign _T_16132 = 6'h6 == _T_10211_60; // @[Mux.scala 46:19:@13136.4]
  assign _T_16133 = _T_16132 ? _T_9260_5 : _T_16131; // @[Mux.scala 46:16:@13137.4]
  assign _T_16134 = 6'h5 == _T_10211_60; // @[Mux.scala 46:19:@13138.4]
  assign _T_16135 = _T_16134 ? _T_9260_4 : _T_16133; // @[Mux.scala 46:16:@13139.4]
  assign _T_16136 = 6'h4 == _T_10211_60; // @[Mux.scala 46:19:@13140.4]
  assign _T_16137 = _T_16136 ? _T_9260_3 : _T_16135; // @[Mux.scala 46:16:@13141.4]
  assign _T_16138 = 6'h3 == _T_10211_60; // @[Mux.scala 46:19:@13142.4]
  assign _T_16139 = _T_16138 ? _T_9260_2 : _T_16137; // @[Mux.scala 46:16:@13143.4]
  assign _T_16140 = 6'h2 == _T_10211_60; // @[Mux.scala 46:19:@13144.4]
  assign _T_16141 = _T_16140 ? _T_9260_1 : _T_16139; // @[Mux.scala 46:16:@13145.4]
  assign _T_16142 = 6'h1 == _T_10211_60; // @[Mux.scala 46:19:@13146.4]
  assign _T_16143 = _T_16142 ? _T_9260_0 : _T_16141; // @[Mux.scala 46:16:@13147.4]
  assign _T_16207 = 6'h3e == _T_10211_61; // @[Mux.scala 46:19:@13149.4]
  assign _T_16208 = _T_16207 ? _T_9260_61 : 8'h0; // @[Mux.scala 46:16:@13150.4]
  assign _T_16209 = 6'h3d == _T_10211_61; // @[Mux.scala 46:19:@13151.4]
  assign _T_16210 = _T_16209 ? _T_9260_60 : _T_16208; // @[Mux.scala 46:16:@13152.4]
  assign _T_16211 = 6'h3c == _T_10211_61; // @[Mux.scala 46:19:@13153.4]
  assign _T_16212 = _T_16211 ? _T_9260_59 : _T_16210; // @[Mux.scala 46:16:@13154.4]
  assign _T_16213 = 6'h3b == _T_10211_61; // @[Mux.scala 46:19:@13155.4]
  assign _T_16214 = _T_16213 ? _T_9260_58 : _T_16212; // @[Mux.scala 46:16:@13156.4]
  assign _T_16215 = 6'h3a == _T_10211_61; // @[Mux.scala 46:19:@13157.4]
  assign _T_16216 = _T_16215 ? _T_9260_57 : _T_16214; // @[Mux.scala 46:16:@13158.4]
  assign _T_16217 = 6'h39 == _T_10211_61; // @[Mux.scala 46:19:@13159.4]
  assign _T_16218 = _T_16217 ? _T_9260_56 : _T_16216; // @[Mux.scala 46:16:@13160.4]
  assign _T_16219 = 6'h38 == _T_10211_61; // @[Mux.scala 46:19:@13161.4]
  assign _T_16220 = _T_16219 ? _T_9260_55 : _T_16218; // @[Mux.scala 46:16:@13162.4]
  assign _T_16221 = 6'h37 == _T_10211_61; // @[Mux.scala 46:19:@13163.4]
  assign _T_16222 = _T_16221 ? _T_9260_54 : _T_16220; // @[Mux.scala 46:16:@13164.4]
  assign _T_16223 = 6'h36 == _T_10211_61; // @[Mux.scala 46:19:@13165.4]
  assign _T_16224 = _T_16223 ? _T_9260_53 : _T_16222; // @[Mux.scala 46:16:@13166.4]
  assign _T_16225 = 6'h35 == _T_10211_61; // @[Mux.scala 46:19:@13167.4]
  assign _T_16226 = _T_16225 ? _T_9260_52 : _T_16224; // @[Mux.scala 46:16:@13168.4]
  assign _T_16227 = 6'h34 == _T_10211_61; // @[Mux.scala 46:19:@13169.4]
  assign _T_16228 = _T_16227 ? _T_9260_51 : _T_16226; // @[Mux.scala 46:16:@13170.4]
  assign _T_16229 = 6'h33 == _T_10211_61; // @[Mux.scala 46:19:@13171.4]
  assign _T_16230 = _T_16229 ? _T_9260_50 : _T_16228; // @[Mux.scala 46:16:@13172.4]
  assign _T_16231 = 6'h32 == _T_10211_61; // @[Mux.scala 46:19:@13173.4]
  assign _T_16232 = _T_16231 ? _T_9260_49 : _T_16230; // @[Mux.scala 46:16:@13174.4]
  assign _T_16233 = 6'h31 == _T_10211_61; // @[Mux.scala 46:19:@13175.4]
  assign _T_16234 = _T_16233 ? _T_9260_48 : _T_16232; // @[Mux.scala 46:16:@13176.4]
  assign _T_16235 = 6'h30 == _T_10211_61; // @[Mux.scala 46:19:@13177.4]
  assign _T_16236 = _T_16235 ? _T_9260_47 : _T_16234; // @[Mux.scala 46:16:@13178.4]
  assign _T_16237 = 6'h2f == _T_10211_61; // @[Mux.scala 46:19:@13179.4]
  assign _T_16238 = _T_16237 ? _T_9260_46 : _T_16236; // @[Mux.scala 46:16:@13180.4]
  assign _T_16239 = 6'h2e == _T_10211_61; // @[Mux.scala 46:19:@13181.4]
  assign _T_16240 = _T_16239 ? _T_9260_45 : _T_16238; // @[Mux.scala 46:16:@13182.4]
  assign _T_16241 = 6'h2d == _T_10211_61; // @[Mux.scala 46:19:@13183.4]
  assign _T_16242 = _T_16241 ? _T_9260_44 : _T_16240; // @[Mux.scala 46:16:@13184.4]
  assign _T_16243 = 6'h2c == _T_10211_61; // @[Mux.scala 46:19:@13185.4]
  assign _T_16244 = _T_16243 ? _T_9260_43 : _T_16242; // @[Mux.scala 46:16:@13186.4]
  assign _T_16245 = 6'h2b == _T_10211_61; // @[Mux.scala 46:19:@13187.4]
  assign _T_16246 = _T_16245 ? _T_9260_42 : _T_16244; // @[Mux.scala 46:16:@13188.4]
  assign _T_16247 = 6'h2a == _T_10211_61; // @[Mux.scala 46:19:@13189.4]
  assign _T_16248 = _T_16247 ? _T_9260_41 : _T_16246; // @[Mux.scala 46:16:@13190.4]
  assign _T_16249 = 6'h29 == _T_10211_61; // @[Mux.scala 46:19:@13191.4]
  assign _T_16250 = _T_16249 ? _T_9260_40 : _T_16248; // @[Mux.scala 46:16:@13192.4]
  assign _T_16251 = 6'h28 == _T_10211_61; // @[Mux.scala 46:19:@13193.4]
  assign _T_16252 = _T_16251 ? _T_9260_39 : _T_16250; // @[Mux.scala 46:16:@13194.4]
  assign _T_16253 = 6'h27 == _T_10211_61; // @[Mux.scala 46:19:@13195.4]
  assign _T_16254 = _T_16253 ? _T_9260_38 : _T_16252; // @[Mux.scala 46:16:@13196.4]
  assign _T_16255 = 6'h26 == _T_10211_61; // @[Mux.scala 46:19:@13197.4]
  assign _T_16256 = _T_16255 ? _T_9260_37 : _T_16254; // @[Mux.scala 46:16:@13198.4]
  assign _T_16257 = 6'h25 == _T_10211_61; // @[Mux.scala 46:19:@13199.4]
  assign _T_16258 = _T_16257 ? _T_9260_36 : _T_16256; // @[Mux.scala 46:16:@13200.4]
  assign _T_16259 = 6'h24 == _T_10211_61; // @[Mux.scala 46:19:@13201.4]
  assign _T_16260 = _T_16259 ? _T_9260_35 : _T_16258; // @[Mux.scala 46:16:@13202.4]
  assign _T_16261 = 6'h23 == _T_10211_61; // @[Mux.scala 46:19:@13203.4]
  assign _T_16262 = _T_16261 ? _T_9260_34 : _T_16260; // @[Mux.scala 46:16:@13204.4]
  assign _T_16263 = 6'h22 == _T_10211_61; // @[Mux.scala 46:19:@13205.4]
  assign _T_16264 = _T_16263 ? _T_9260_33 : _T_16262; // @[Mux.scala 46:16:@13206.4]
  assign _T_16265 = 6'h21 == _T_10211_61; // @[Mux.scala 46:19:@13207.4]
  assign _T_16266 = _T_16265 ? _T_9260_32 : _T_16264; // @[Mux.scala 46:16:@13208.4]
  assign _T_16267 = 6'h20 == _T_10211_61; // @[Mux.scala 46:19:@13209.4]
  assign _T_16268 = _T_16267 ? _T_9260_31 : _T_16266; // @[Mux.scala 46:16:@13210.4]
  assign _T_16269 = 6'h1f == _T_10211_61; // @[Mux.scala 46:19:@13211.4]
  assign _T_16270 = _T_16269 ? _T_9260_30 : _T_16268; // @[Mux.scala 46:16:@13212.4]
  assign _T_16271 = 6'h1e == _T_10211_61; // @[Mux.scala 46:19:@13213.4]
  assign _T_16272 = _T_16271 ? _T_9260_29 : _T_16270; // @[Mux.scala 46:16:@13214.4]
  assign _T_16273 = 6'h1d == _T_10211_61; // @[Mux.scala 46:19:@13215.4]
  assign _T_16274 = _T_16273 ? _T_9260_28 : _T_16272; // @[Mux.scala 46:16:@13216.4]
  assign _T_16275 = 6'h1c == _T_10211_61; // @[Mux.scala 46:19:@13217.4]
  assign _T_16276 = _T_16275 ? _T_9260_27 : _T_16274; // @[Mux.scala 46:16:@13218.4]
  assign _T_16277 = 6'h1b == _T_10211_61; // @[Mux.scala 46:19:@13219.4]
  assign _T_16278 = _T_16277 ? _T_9260_26 : _T_16276; // @[Mux.scala 46:16:@13220.4]
  assign _T_16279 = 6'h1a == _T_10211_61; // @[Mux.scala 46:19:@13221.4]
  assign _T_16280 = _T_16279 ? _T_9260_25 : _T_16278; // @[Mux.scala 46:16:@13222.4]
  assign _T_16281 = 6'h19 == _T_10211_61; // @[Mux.scala 46:19:@13223.4]
  assign _T_16282 = _T_16281 ? _T_9260_24 : _T_16280; // @[Mux.scala 46:16:@13224.4]
  assign _T_16283 = 6'h18 == _T_10211_61; // @[Mux.scala 46:19:@13225.4]
  assign _T_16284 = _T_16283 ? _T_9260_23 : _T_16282; // @[Mux.scala 46:16:@13226.4]
  assign _T_16285 = 6'h17 == _T_10211_61; // @[Mux.scala 46:19:@13227.4]
  assign _T_16286 = _T_16285 ? _T_9260_22 : _T_16284; // @[Mux.scala 46:16:@13228.4]
  assign _T_16287 = 6'h16 == _T_10211_61; // @[Mux.scala 46:19:@13229.4]
  assign _T_16288 = _T_16287 ? _T_9260_21 : _T_16286; // @[Mux.scala 46:16:@13230.4]
  assign _T_16289 = 6'h15 == _T_10211_61; // @[Mux.scala 46:19:@13231.4]
  assign _T_16290 = _T_16289 ? _T_9260_20 : _T_16288; // @[Mux.scala 46:16:@13232.4]
  assign _T_16291 = 6'h14 == _T_10211_61; // @[Mux.scala 46:19:@13233.4]
  assign _T_16292 = _T_16291 ? _T_9260_19 : _T_16290; // @[Mux.scala 46:16:@13234.4]
  assign _T_16293 = 6'h13 == _T_10211_61; // @[Mux.scala 46:19:@13235.4]
  assign _T_16294 = _T_16293 ? _T_9260_18 : _T_16292; // @[Mux.scala 46:16:@13236.4]
  assign _T_16295 = 6'h12 == _T_10211_61; // @[Mux.scala 46:19:@13237.4]
  assign _T_16296 = _T_16295 ? _T_9260_17 : _T_16294; // @[Mux.scala 46:16:@13238.4]
  assign _T_16297 = 6'h11 == _T_10211_61; // @[Mux.scala 46:19:@13239.4]
  assign _T_16298 = _T_16297 ? _T_9260_16 : _T_16296; // @[Mux.scala 46:16:@13240.4]
  assign _T_16299 = 6'h10 == _T_10211_61; // @[Mux.scala 46:19:@13241.4]
  assign _T_16300 = _T_16299 ? _T_9260_15 : _T_16298; // @[Mux.scala 46:16:@13242.4]
  assign _T_16301 = 6'hf == _T_10211_61; // @[Mux.scala 46:19:@13243.4]
  assign _T_16302 = _T_16301 ? _T_9260_14 : _T_16300; // @[Mux.scala 46:16:@13244.4]
  assign _T_16303 = 6'he == _T_10211_61; // @[Mux.scala 46:19:@13245.4]
  assign _T_16304 = _T_16303 ? _T_9260_13 : _T_16302; // @[Mux.scala 46:16:@13246.4]
  assign _T_16305 = 6'hd == _T_10211_61; // @[Mux.scala 46:19:@13247.4]
  assign _T_16306 = _T_16305 ? _T_9260_12 : _T_16304; // @[Mux.scala 46:16:@13248.4]
  assign _T_16307 = 6'hc == _T_10211_61; // @[Mux.scala 46:19:@13249.4]
  assign _T_16308 = _T_16307 ? _T_9260_11 : _T_16306; // @[Mux.scala 46:16:@13250.4]
  assign _T_16309 = 6'hb == _T_10211_61; // @[Mux.scala 46:19:@13251.4]
  assign _T_16310 = _T_16309 ? _T_9260_10 : _T_16308; // @[Mux.scala 46:16:@13252.4]
  assign _T_16311 = 6'ha == _T_10211_61; // @[Mux.scala 46:19:@13253.4]
  assign _T_16312 = _T_16311 ? _T_9260_9 : _T_16310; // @[Mux.scala 46:16:@13254.4]
  assign _T_16313 = 6'h9 == _T_10211_61; // @[Mux.scala 46:19:@13255.4]
  assign _T_16314 = _T_16313 ? _T_9260_8 : _T_16312; // @[Mux.scala 46:16:@13256.4]
  assign _T_16315 = 6'h8 == _T_10211_61; // @[Mux.scala 46:19:@13257.4]
  assign _T_16316 = _T_16315 ? _T_9260_7 : _T_16314; // @[Mux.scala 46:16:@13258.4]
  assign _T_16317 = 6'h7 == _T_10211_61; // @[Mux.scala 46:19:@13259.4]
  assign _T_16318 = _T_16317 ? _T_9260_6 : _T_16316; // @[Mux.scala 46:16:@13260.4]
  assign _T_16319 = 6'h6 == _T_10211_61; // @[Mux.scala 46:19:@13261.4]
  assign _T_16320 = _T_16319 ? _T_9260_5 : _T_16318; // @[Mux.scala 46:16:@13262.4]
  assign _T_16321 = 6'h5 == _T_10211_61; // @[Mux.scala 46:19:@13263.4]
  assign _T_16322 = _T_16321 ? _T_9260_4 : _T_16320; // @[Mux.scala 46:16:@13264.4]
  assign _T_16323 = 6'h4 == _T_10211_61; // @[Mux.scala 46:19:@13265.4]
  assign _T_16324 = _T_16323 ? _T_9260_3 : _T_16322; // @[Mux.scala 46:16:@13266.4]
  assign _T_16325 = 6'h3 == _T_10211_61; // @[Mux.scala 46:19:@13267.4]
  assign _T_16326 = _T_16325 ? _T_9260_2 : _T_16324; // @[Mux.scala 46:16:@13268.4]
  assign _T_16327 = 6'h2 == _T_10211_61; // @[Mux.scala 46:19:@13269.4]
  assign _T_16328 = _T_16327 ? _T_9260_1 : _T_16326; // @[Mux.scala 46:16:@13270.4]
  assign _T_16329 = 6'h1 == _T_10211_61; // @[Mux.scala 46:19:@13271.4]
  assign _T_16330 = _T_16329 ? _T_9260_0 : _T_16328; // @[Mux.scala 46:16:@13272.4]
  assign _T_16395 = 6'h3f == _T_10211_62; // @[Mux.scala 46:19:@13274.4]
  assign _T_16396 = _T_16395 ? _T_9260_62 : 8'h0; // @[Mux.scala 46:16:@13275.4]
  assign _T_16397 = 6'h3e == _T_10211_62; // @[Mux.scala 46:19:@13276.4]
  assign _T_16398 = _T_16397 ? _T_9260_61 : _T_16396; // @[Mux.scala 46:16:@13277.4]
  assign _T_16399 = 6'h3d == _T_10211_62; // @[Mux.scala 46:19:@13278.4]
  assign _T_16400 = _T_16399 ? _T_9260_60 : _T_16398; // @[Mux.scala 46:16:@13279.4]
  assign _T_16401 = 6'h3c == _T_10211_62; // @[Mux.scala 46:19:@13280.4]
  assign _T_16402 = _T_16401 ? _T_9260_59 : _T_16400; // @[Mux.scala 46:16:@13281.4]
  assign _T_16403 = 6'h3b == _T_10211_62; // @[Mux.scala 46:19:@13282.4]
  assign _T_16404 = _T_16403 ? _T_9260_58 : _T_16402; // @[Mux.scala 46:16:@13283.4]
  assign _T_16405 = 6'h3a == _T_10211_62; // @[Mux.scala 46:19:@13284.4]
  assign _T_16406 = _T_16405 ? _T_9260_57 : _T_16404; // @[Mux.scala 46:16:@13285.4]
  assign _T_16407 = 6'h39 == _T_10211_62; // @[Mux.scala 46:19:@13286.4]
  assign _T_16408 = _T_16407 ? _T_9260_56 : _T_16406; // @[Mux.scala 46:16:@13287.4]
  assign _T_16409 = 6'h38 == _T_10211_62; // @[Mux.scala 46:19:@13288.4]
  assign _T_16410 = _T_16409 ? _T_9260_55 : _T_16408; // @[Mux.scala 46:16:@13289.4]
  assign _T_16411 = 6'h37 == _T_10211_62; // @[Mux.scala 46:19:@13290.4]
  assign _T_16412 = _T_16411 ? _T_9260_54 : _T_16410; // @[Mux.scala 46:16:@13291.4]
  assign _T_16413 = 6'h36 == _T_10211_62; // @[Mux.scala 46:19:@13292.4]
  assign _T_16414 = _T_16413 ? _T_9260_53 : _T_16412; // @[Mux.scala 46:16:@13293.4]
  assign _T_16415 = 6'h35 == _T_10211_62; // @[Mux.scala 46:19:@13294.4]
  assign _T_16416 = _T_16415 ? _T_9260_52 : _T_16414; // @[Mux.scala 46:16:@13295.4]
  assign _T_16417 = 6'h34 == _T_10211_62; // @[Mux.scala 46:19:@13296.4]
  assign _T_16418 = _T_16417 ? _T_9260_51 : _T_16416; // @[Mux.scala 46:16:@13297.4]
  assign _T_16419 = 6'h33 == _T_10211_62; // @[Mux.scala 46:19:@13298.4]
  assign _T_16420 = _T_16419 ? _T_9260_50 : _T_16418; // @[Mux.scala 46:16:@13299.4]
  assign _T_16421 = 6'h32 == _T_10211_62; // @[Mux.scala 46:19:@13300.4]
  assign _T_16422 = _T_16421 ? _T_9260_49 : _T_16420; // @[Mux.scala 46:16:@13301.4]
  assign _T_16423 = 6'h31 == _T_10211_62; // @[Mux.scala 46:19:@13302.4]
  assign _T_16424 = _T_16423 ? _T_9260_48 : _T_16422; // @[Mux.scala 46:16:@13303.4]
  assign _T_16425 = 6'h30 == _T_10211_62; // @[Mux.scala 46:19:@13304.4]
  assign _T_16426 = _T_16425 ? _T_9260_47 : _T_16424; // @[Mux.scala 46:16:@13305.4]
  assign _T_16427 = 6'h2f == _T_10211_62; // @[Mux.scala 46:19:@13306.4]
  assign _T_16428 = _T_16427 ? _T_9260_46 : _T_16426; // @[Mux.scala 46:16:@13307.4]
  assign _T_16429 = 6'h2e == _T_10211_62; // @[Mux.scala 46:19:@13308.4]
  assign _T_16430 = _T_16429 ? _T_9260_45 : _T_16428; // @[Mux.scala 46:16:@13309.4]
  assign _T_16431 = 6'h2d == _T_10211_62; // @[Mux.scala 46:19:@13310.4]
  assign _T_16432 = _T_16431 ? _T_9260_44 : _T_16430; // @[Mux.scala 46:16:@13311.4]
  assign _T_16433 = 6'h2c == _T_10211_62; // @[Mux.scala 46:19:@13312.4]
  assign _T_16434 = _T_16433 ? _T_9260_43 : _T_16432; // @[Mux.scala 46:16:@13313.4]
  assign _T_16435 = 6'h2b == _T_10211_62; // @[Mux.scala 46:19:@13314.4]
  assign _T_16436 = _T_16435 ? _T_9260_42 : _T_16434; // @[Mux.scala 46:16:@13315.4]
  assign _T_16437 = 6'h2a == _T_10211_62; // @[Mux.scala 46:19:@13316.4]
  assign _T_16438 = _T_16437 ? _T_9260_41 : _T_16436; // @[Mux.scala 46:16:@13317.4]
  assign _T_16439 = 6'h29 == _T_10211_62; // @[Mux.scala 46:19:@13318.4]
  assign _T_16440 = _T_16439 ? _T_9260_40 : _T_16438; // @[Mux.scala 46:16:@13319.4]
  assign _T_16441 = 6'h28 == _T_10211_62; // @[Mux.scala 46:19:@13320.4]
  assign _T_16442 = _T_16441 ? _T_9260_39 : _T_16440; // @[Mux.scala 46:16:@13321.4]
  assign _T_16443 = 6'h27 == _T_10211_62; // @[Mux.scala 46:19:@13322.4]
  assign _T_16444 = _T_16443 ? _T_9260_38 : _T_16442; // @[Mux.scala 46:16:@13323.4]
  assign _T_16445 = 6'h26 == _T_10211_62; // @[Mux.scala 46:19:@13324.4]
  assign _T_16446 = _T_16445 ? _T_9260_37 : _T_16444; // @[Mux.scala 46:16:@13325.4]
  assign _T_16447 = 6'h25 == _T_10211_62; // @[Mux.scala 46:19:@13326.4]
  assign _T_16448 = _T_16447 ? _T_9260_36 : _T_16446; // @[Mux.scala 46:16:@13327.4]
  assign _T_16449 = 6'h24 == _T_10211_62; // @[Mux.scala 46:19:@13328.4]
  assign _T_16450 = _T_16449 ? _T_9260_35 : _T_16448; // @[Mux.scala 46:16:@13329.4]
  assign _T_16451 = 6'h23 == _T_10211_62; // @[Mux.scala 46:19:@13330.4]
  assign _T_16452 = _T_16451 ? _T_9260_34 : _T_16450; // @[Mux.scala 46:16:@13331.4]
  assign _T_16453 = 6'h22 == _T_10211_62; // @[Mux.scala 46:19:@13332.4]
  assign _T_16454 = _T_16453 ? _T_9260_33 : _T_16452; // @[Mux.scala 46:16:@13333.4]
  assign _T_16455 = 6'h21 == _T_10211_62; // @[Mux.scala 46:19:@13334.4]
  assign _T_16456 = _T_16455 ? _T_9260_32 : _T_16454; // @[Mux.scala 46:16:@13335.4]
  assign _T_16457 = 6'h20 == _T_10211_62; // @[Mux.scala 46:19:@13336.4]
  assign _T_16458 = _T_16457 ? _T_9260_31 : _T_16456; // @[Mux.scala 46:16:@13337.4]
  assign _T_16459 = 6'h1f == _T_10211_62; // @[Mux.scala 46:19:@13338.4]
  assign _T_16460 = _T_16459 ? _T_9260_30 : _T_16458; // @[Mux.scala 46:16:@13339.4]
  assign _T_16461 = 6'h1e == _T_10211_62; // @[Mux.scala 46:19:@13340.4]
  assign _T_16462 = _T_16461 ? _T_9260_29 : _T_16460; // @[Mux.scala 46:16:@13341.4]
  assign _T_16463 = 6'h1d == _T_10211_62; // @[Mux.scala 46:19:@13342.4]
  assign _T_16464 = _T_16463 ? _T_9260_28 : _T_16462; // @[Mux.scala 46:16:@13343.4]
  assign _T_16465 = 6'h1c == _T_10211_62; // @[Mux.scala 46:19:@13344.4]
  assign _T_16466 = _T_16465 ? _T_9260_27 : _T_16464; // @[Mux.scala 46:16:@13345.4]
  assign _T_16467 = 6'h1b == _T_10211_62; // @[Mux.scala 46:19:@13346.4]
  assign _T_16468 = _T_16467 ? _T_9260_26 : _T_16466; // @[Mux.scala 46:16:@13347.4]
  assign _T_16469 = 6'h1a == _T_10211_62; // @[Mux.scala 46:19:@13348.4]
  assign _T_16470 = _T_16469 ? _T_9260_25 : _T_16468; // @[Mux.scala 46:16:@13349.4]
  assign _T_16471 = 6'h19 == _T_10211_62; // @[Mux.scala 46:19:@13350.4]
  assign _T_16472 = _T_16471 ? _T_9260_24 : _T_16470; // @[Mux.scala 46:16:@13351.4]
  assign _T_16473 = 6'h18 == _T_10211_62; // @[Mux.scala 46:19:@13352.4]
  assign _T_16474 = _T_16473 ? _T_9260_23 : _T_16472; // @[Mux.scala 46:16:@13353.4]
  assign _T_16475 = 6'h17 == _T_10211_62; // @[Mux.scala 46:19:@13354.4]
  assign _T_16476 = _T_16475 ? _T_9260_22 : _T_16474; // @[Mux.scala 46:16:@13355.4]
  assign _T_16477 = 6'h16 == _T_10211_62; // @[Mux.scala 46:19:@13356.4]
  assign _T_16478 = _T_16477 ? _T_9260_21 : _T_16476; // @[Mux.scala 46:16:@13357.4]
  assign _T_16479 = 6'h15 == _T_10211_62; // @[Mux.scala 46:19:@13358.4]
  assign _T_16480 = _T_16479 ? _T_9260_20 : _T_16478; // @[Mux.scala 46:16:@13359.4]
  assign _T_16481 = 6'h14 == _T_10211_62; // @[Mux.scala 46:19:@13360.4]
  assign _T_16482 = _T_16481 ? _T_9260_19 : _T_16480; // @[Mux.scala 46:16:@13361.4]
  assign _T_16483 = 6'h13 == _T_10211_62; // @[Mux.scala 46:19:@13362.4]
  assign _T_16484 = _T_16483 ? _T_9260_18 : _T_16482; // @[Mux.scala 46:16:@13363.4]
  assign _T_16485 = 6'h12 == _T_10211_62; // @[Mux.scala 46:19:@13364.4]
  assign _T_16486 = _T_16485 ? _T_9260_17 : _T_16484; // @[Mux.scala 46:16:@13365.4]
  assign _T_16487 = 6'h11 == _T_10211_62; // @[Mux.scala 46:19:@13366.4]
  assign _T_16488 = _T_16487 ? _T_9260_16 : _T_16486; // @[Mux.scala 46:16:@13367.4]
  assign _T_16489 = 6'h10 == _T_10211_62; // @[Mux.scala 46:19:@13368.4]
  assign _T_16490 = _T_16489 ? _T_9260_15 : _T_16488; // @[Mux.scala 46:16:@13369.4]
  assign _T_16491 = 6'hf == _T_10211_62; // @[Mux.scala 46:19:@13370.4]
  assign _T_16492 = _T_16491 ? _T_9260_14 : _T_16490; // @[Mux.scala 46:16:@13371.4]
  assign _T_16493 = 6'he == _T_10211_62; // @[Mux.scala 46:19:@13372.4]
  assign _T_16494 = _T_16493 ? _T_9260_13 : _T_16492; // @[Mux.scala 46:16:@13373.4]
  assign _T_16495 = 6'hd == _T_10211_62; // @[Mux.scala 46:19:@13374.4]
  assign _T_16496 = _T_16495 ? _T_9260_12 : _T_16494; // @[Mux.scala 46:16:@13375.4]
  assign _T_16497 = 6'hc == _T_10211_62; // @[Mux.scala 46:19:@13376.4]
  assign _T_16498 = _T_16497 ? _T_9260_11 : _T_16496; // @[Mux.scala 46:16:@13377.4]
  assign _T_16499 = 6'hb == _T_10211_62; // @[Mux.scala 46:19:@13378.4]
  assign _T_16500 = _T_16499 ? _T_9260_10 : _T_16498; // @[Mux.scala 46:16:@13379.4]
  assign _T_16501 = 6'ha == _T_10211_62; // @[Mux.scala 46:19:@13380.4]
  assign _T_16502 = _T_16501 ? _T_9260_9 : _T_16500; // @[Mux.scala 46:16:@13381.4]
  assign _T_16503 = 6'h9 == _T_10211_62; // @[Mux.scala 46:19:@13382.4]
  assign _T_16504 = _T_16503 ? _T_9260_8 : _T_16502; // @[Mux.scala 46:16:@13383.4]
  assign _T_16505 = 6'h8 == _T_10211_62; // @[Mux.scala 46:19:@13384.4]
  assign _T_16506 = _T_16505 ? _T_9260_7 : _T_16504; // @[Mux.scala 46:16:@13385.4]
  assign _T_16507 = 6'h7 == _T_10211_62; // @[Mux.scala 46:19:@13386.4]
  assign _T_16508 = _T_16507 ? _T_9260_6 : _T_16506; // @[Mux.scala 46:16:@13387.4]
  assign _T_16509 = 6'h6 == _T_10211_62; // @[Mux.scala 46:19:@13388.4]
  assign _T_16510 = _T_16509 ? _T_9260_5 : _T_16508; // @[Mux.scala 46:16:@13389.4]
  assign _T_16511 = 6'h5 == _T_10211_62; // @[Mux.scala 46:19:@13390.4]
  assign _T_16512 = _T_16511 ? _T_9260_4 : _T_16510; // @[Mux.scala 46:16:@13391.4]
  assign _T_16513 = 6'h4 == _T_10211_62; // @[Mux.scala 46:19:@13392.4]
  assign _T_16514 = _T_16513 ? _T_9260_3 : _T_16512; // @[Mux.scala 46:16:@13393.4]
  assign _T_16515 = 6'h3 == _T_10211_62; // @[Mux.scala 46:19:@13394.4]
  assign _T_16516 = _T_16515 ? _T_9260_2 : _T_16514; // @[Mux.scala 46:16:@13395.4]
  assign _T_16517 = 6'h2 == _T_10211_62; // @[Mux.scala 46:19:@13396.4]
  assign _T_16518 = _T_16517 ? _T_9260_1 : _T_16516; // @[Mux.scala 46:16:@13397.4]
  assign _T_16519 = 6'h1 == _T_10211_62; // @[Mux.scala 46:19:@13398.4]
  assign _T_16520 = _T_16519 ? _T_9260_0 : _T_16518; // @[Mux.scala 46:16:@13399.4]
  assign _T_16586 = 7'h40 == _T_10211_63; // @[Mux.scala 46:19:@13401.4]
  assign _T_16587 = _T_16586 ? _T_9260_63 : 8'h0; // @[Mux.scala 46:16:@13402.4]
  assign _T_16588 = 7'h3f == _T_10211_63; // @[Mux.scala 46:19:@13403.4]
  assign _T_16589 = _T_16588 ? _T_9260_62 : _T_16587; // @[Mux.scala 46:16:@13404.4]
  assign _T_16590 = 7'h3e == _T_10211_63; // @[Mux.scala 46:19:@13405.4]
  assign _T_16591 = _T_16590 ? _T_9260_61 : _T_16589; // @[Mux.scala 46:16:@13406.4]
  assign _T_16592 = 7'h3d == _T_10211_63; // @[Mux.scala 46:19:@13407.4]
  assign _T_16593 = _T_16592 ? _T_9260_60 : _T_16591; // @[Mux.scala 46:16:@13408.4]
  assign _T_16594 = 7'h3c == _T_10211_63; // @[Mux.scala 46:19:@13409.4]
  assign _T_16595 = _T_16594 ? _T_9260_59 : _T_16593; // @[Mux.scala 46:16:@13410.4]
  assign _T_16596 = 7'h3b == _T_10211_63; // @[Mux.scala 46:19:@13411.4]
  assign _T_16597 = _T_16596 ? _T_9260_58 : _T_16595; // @[Mux.scala 46:16:@13412.4]
  assign _T_16598 = 7'h3a == _T_10211_63; // @[Mux.scala 46:19:@13413.4]
  assign _T_16599 = _T_16598 ? _T_9260_57 : _T_16597; // @[Mux.scala 46:16:@13414.4]
  assign _T_16600 = 7'h39 == _T_10211_63; // @[Mux.scala 46:19:@13415.4]
  assign _T_16601 = _T_16600 ? _T_9260_56 : _T_16599; // @[Mux.scala 46:16:@13416.4]
  assign _T_16602 = 7'h38 == _T_10211_63; // @[Mux.scala 46:19:@13417.4]
  assign _T_16603 = _T_16602 ? _T_9260_55 : _T_16601; // @[Mux.scala 46:16:@13418.4]
  assign _T_16604 = 7'h37 == _T_10211_63; // @[Mux.scala 46:19:@13419.4]
  assign _T_16605 = _T_16604 ? _T_9260_54 : _T_16603; // @[Mux.scala 46:16:@13420.4]
  assign _T_16606 = 7'h36 == _T_10211_63; // @[Mux.scala 46:19:@13421.4]
  assign _T_16607 = _T_16606 ? _T_9260_53 : _T_16605; // @[Mux.scala 46:16:@13422.4]
  assign _T_16608 = 7'h35 == _T_10211_63; // @[Mux.scala 46:19:@13423.4]
  assign _T_16609 = _T_16608 ? _T_9260_52 : _T_16607; // @[Mux.scala 46:16:@13424.4]
  assign _T_16610 = 7'h34 == _T_10211_63; // @[Mux.scala 46:19:@13425.4]
  assign _T_16611 = _T_16610 ? _T_9260_51 : _T_16609; // @[Mux.scala 46:16:@13426.4]
  assign _T_16612 = 7'h33 == _T_10211_63; // @[Mux.scala 46:19:@13427.4]
  assign _T_16613 = _T_16612 ? _T_9260_50 : _T_16611; // @[Mux.scala 46:16:@13428.4]
  assign _T_16614 = 7'h32 == _T_10211_63; // @[Mux.scala 46:19:@13429.4]
  assign _T_16615 = _T_16614 ? _T_9260_49 : _T_16613; // @[Mux.scala 46:16:@13430.4]
  assign _T_16616 = 7'h31 == _T_10211_63; // @[Mux.scala 46:19:@13431.4]
  assign _T_16617 = _T_16616 ? _T_9260_48 : _T_16615; // @[Mux.scala 46:16:@13432.4]
  assign _T_16618 = 7'h30 == _T_10211_63; // @[Mux.scala 46:19:@13433.4]
  assign _T_16619 = _T_16618 ? _T_9260_47 : _T_16617; // @[Mux.scala 46:16:@13434.4]
  assign _T_16620 = 7'h2f == _T_10211_63; // @[Mux.scala 46:19:@13435.4]
  assign _T_16621 = _T_16620 ? _T_9260_46 : _T_16619; // @[Mux.scala 46:16:@13436.4]
  assign _T_16622 = 7'h2e == _T_10211_63; // @[Mux.scala 46:19:@13437.4]
  assign _T_16623 = _T_16622 ? _T_9260_45 : _T_16621; // @[Mux.scala 46:16:@13438.4]
  assign _T_16624 = 7'h2d == _T_10211_63; // @[Mux.scala 46:19:@13439.4]
  assign _T_16625 = _T_16624 ? _T_9260_44 : _T_16623; // @[Mux.scala 46:16:@13440.4]
  assign _T_16626 = 7'h2c == _T_10211_63; // @[Mux.scala 46:19:@13441.4]
  assign _T_16627 = _T_16626 ? _T_9260_43 : _T_16625; // @[Mux.scala 46:16:@13442.4]
  assign _T_16628 = 7'h2b == _T_10211_63; // @[Mux.scala 46:19:@13443.4]
  assign _T_16629 = _T_16628 ? _T_9260_42 : _T_16627; // @[Mux.scala 46:16:@13444.4]
  assign _T_16630 = 7'h2a == _T_10211_63; // @[Mux.scala 46:19:@13445.4]
  assign _T_16631 = _T_16630 ? _T_9260_41 : _T_16629; // @[Mux.scala 46:16:@13446.4]
  assign _T_16632 = 7'h29 == _T_10211_63; // @[Mux.scala 46:19:@13447.4]
  assign _T_16633 = _T_16632 ? _T_9260_40 : _T_16631; // @[Mux.scala 46:16:@13448.4]
  assign _T_16634 = 7'h28 == _T_10211_63; // @[Mux.scala 46:19:@13449.4]
  assign _T_16635 = _T_16634 ? _T_9260_39 : _T_16633; // @[Mux.scala 46:16:@13450.4]
  assign _T_16636 = 7'h27 == _T_10211_63; // @[Mux.scala 46:19:@13451.4]
  assign _T_16637 = _T_16636 ? _T_9260_38 : _T_16635; // @[Mux.scala 46:16:@13452.4]
  assign _T_16638 = 7'h26 == _T_10211_63; // @[Mux.scala 46:19:@13453.4]
  assign _T_16639 = _T_16638 ? _T_9260_37 : _T_16637; // @[Mux.scala 46:16:@13454.4]
  assign _T_16640 = 7'h25 == _T_10211_63; // @[Mux.scala 46:19:@13455.4]
  assign _T_16641 = _T_16640 ? _T_9260_36 : _T_16639; // @[Mux.scala 46:16:@13456.4]
  assign _T_16642 = 7'h24 == _T_10211_63; // @[Mux.scala 46:19:@13457.4]
  assign _T_16643 = _T_16642 ? _T_9260_35 : _T_16641; // @[Mux.scala 46:16:@13458.4]
  assign _T_16644 = 7'h23 == _T_10211_63; // @[Mux.scala 46:19:@13459.4]
  assign _T_16645 = _T_16644 ? _T_9260_34 : _T_16643; // @[Mux.scala 46:16:@13460.4]
  assign _T_16646 = 7'h22 == _T_10211_63; // @[Mux.scala 46:19:@13461.4]
  assign _T_16647 = _T_16646 ? _T_9260_33 : _T_16645; // @[Mux.scala 46:16:@13462.4]
  assign _T_16648 = 7'h21 == _T_10211_63; // @[Mux.scala 46:19:@13463.4]
  assign _T_16649 = _T_16648 ? _T_9260_32 : _T_16647; // @[Mux.scala 46:16:@13464.4]
  assign _T_16650 = 7'h20 == _T_10211_63; // @[Mux.scala 46:19:@13465.4]
  assign _T_16651 = _T_16650 ? _T_9260_31 : _T_16649; // @[Mux.scala 46:16:@13466.4]
  assign _T_16652 = 7'h1f == _T_10211_63; // @[Mux.scala 46:19:@13467.4]
  assign _T_16653 = _T_16652 ? _T_9260_30 : _T_16651; // @[Mux.scala 46:16:@13468.4]
  assign _T_16654 = 7'h1e == _T_10211_63; // @[Mux.scala 46:19:@13469.4]
  assign _T_16655 = _T_16654 ? _T_9260_29 : _T_16653; // @[Mux.scala 46:16:@13470.4]
  assign _T_16656 = 7'h1d == _T_10211_63; // @[Mux.scala 46:19:@13471.4]
  assign _T_16657 = _T_16656 ? _T_9260_28 : _T_16655; // @[Mux.scala 46:16:@13472.4]
  assign _T_16658 = 7'h1c == _T_10211_63; // @[Mux.scala 46:19:@13473.4]
  assign _T_16659 = _T_16658 ? _T_9260_27 : _T_16657; // @[Mux.scala 46:16:@13474.4]
  assign _T_16660 = 7'h1b == _T_10211_63; // @[Mux.scala 46:19:@13475.4]
  assign _T_16661 = _T_16660 ? _T_9260_26 : _T_16659; // @[Mux.scala 46:16:@13476.4]
  assign _T_16662 = 7'h1a == _T_10211_63; // @[Mux.scala 46:19:@13477.4]
  assign _T_16663 = _T_16662 ? _T_9260_25 : _T_16661; // @[Mux.scala 46:16:@13478.4]
  assign _T_16664 = 7'h19 == _T_10211_63; // @[Mux.scala 46:19:@13479.4]
  assign _T_16665 = _T_16664 ? _T_9260_24 : _T_16663; // @[Mux.scala 46:16:@13480.4]
  assign _T_16666 = 7'h18 == _T_10211_63; // @[Mux.scala 46:19:@13481.4]
  assign _T_16667 = _T_16666 ? _T_9260_23 : _T_16665; // @[Mux.scala 46:16:@13482.4]
  assign _T_16668 = 7'h17 == _T_10211_63; // @[Mux.scala 46:19:@13483.4]
  assign _T_16669 = _T_16668 ? _T_9260_22 : _T_16667; // @[Mux.scala 46:16:@13484.4]
  assign _T_16670 = 7'h16 == _T_10211_63; // @[Mux.scala 46:19:@13485.4]
  assign _T_16671 = _T_16670 ? _T_9260_21 : _T_16669; // @[Mux.scala 46:16:@13486.4]
  assign _T_16672 = 7'h15 == _T_10211_63; // @[Mux.scala 46:19:@13487.4]
  assign _T_16673 = _T_16672 ? _T_9260_20 : _T_16671; // @[Mux.scala 46:16:@13488.4]
  assign _T_16674 = 7'h14 == _T_10211_63; // @[Mux.scala 46:19:@13489.4]
  assign _T_16675 = _T_16674 ? _T_9260_19 : _T_16673; // @[Mux.scala 46:16:@13490.4]
  assign _T_16676 = 7'h13 == _T_10211_63; // @[Mux.scala 46:19:@13491.4]
  assign _T_16677 = _T_16676 ? _T_9260_18 : _T_16675; // @[Mux.scala 46:16:@13492.4]
  assign _T_16678 = 7'h12 == _T_10211_63; // @[Mux.scala 46:19:@13493.4]
  assign _T_16679 = _T_16678 ? _T_9260_17 : _T_16677; // @[Mux.scala 46:16:@13494.4]
  assign _T_16680 = 7'h11 == _T_10211_63; // @[Mux.scala 46:19:@13495.4]
  assign _T_16681 = _T_16680 ? _T_9260_16 : _T_16679; // @[Mux.scala 46:16:@13496.4]
  assign _T_16682 = 7'h10 == _T_10211_63; // @[Mux.scala 46:19:@13497.4]
  assign _T_16683 = _T_16682 ? _T_9260_15 : _T_16681; // @[Mux.scala 46:16:@13498.4]
  assign _T_16684 = 7'hf == _T_10211_63; // @[Mux.scala 46:19:@13499.4]
  assign _T_16685 = _T_16684 ? _T_9260_14 : _T_16683; // @[Mux.scala 46:16:@13500.4]
  assign _T_16686 = 7'he == _T_10211_63; // @[Mux.scala 46:19:@13501.4]
  assign _T_16687 = _T_16686 ? _T_9260_13 : _T_16685; // @[Mux.scala 46:16:@13502.4]
  assign _T_16688 = 7'hd == _T_10211_63; // @[Mux.scala 46:19:@13503.4]
  assign _T_16689 = _T_16688 ? _T_9260_12 : _T_16687; // @[Mux.scala 46:16:@13504.4]
  assign _T_16690 = 7'hc == _T_10211_63; // @[Mux.scala 46:19:@13505.4]
  assign _T_16691 = _T_16690 ? _T_9260_11 : _T_16689; // @[Mux.scala 46:16:@13506.4]
  assign _T_16692 = 7'hb == _T_10211_63; // @[Mux.scala 46:19:@13507.4]
  assign _T_16693 = _T_16692 ? _T_9260_10 : _T_16691; // @[Mux.scala 46:16:@13508.4]
  assign _T_16694 = 7'ha == _T_10211_63; // @[Mux.scala 46:19:@13509.4]
  assign _T_16695 = _T_16694 ? _T_9260_9 : _T_16693; // @[Mux.scala 46:16:@13510.4]
  assign _T_16696 = 7'h9 == _T_10211_63; // @[Mux.scala 46:19:@13511.4]
  assign _T_16697 = _T_16696 ? _T_9260_8 : _T_16695; // @[Mux.scala 46:16:@13512.4]
  assign _T_16698 = 7'h8 == _T_10211_63; // @[Mux.scala 46:19:@13513.4]
  assign _T_16699 = _T_16698 ? _T_9260_7 : _T_16697; // @[Mux.scala 46:16:@13514.4]
  assign _T_16700 = 7'h7 == _T_10211_63; // @[Mux.scala 46:19:@13515.4]
  assign _T_16701 = _T_16700 ? _T_9260_6 : _T_16699; // @[Mux.scala 46:16:@13516.4]
  assign _T_16702 = 7'h6 == _T_10211_63; // @[Mux.scala 46:19:@13517.4]
  assign _T_16703 = _T_16702 ? _T_9260_5 : _T_16701; // @[Mux.scala 46:16:@13518.4]
  assign _T_16704 = 7'h5 == _T_10211_63; // @[Mux.scala 46:19:@13519.4]
  assign _T_16705 = _T_16704 ? _T_9260_4 : _T_16703; // @[Mux.scala 46:16:@13520.4]
  assign _T_16706 = 7'h4 == _T_10211_63; // @[Mux.scala 46:19:@13521.4]
  assign _T_16707 = _T_16706 ? _T_9260_3 : _T_16705; // @[Mux.scala 46:16:@13522.4]
  assign _T_16708 = 7'h3 == _T_10211_63; // @[Mux.scala 46:19:@13523.4]
  assign _T_16709 = _T_16708 ? _T_9260_2 : _T_16707; // @[Mux.scala 46:16:@13524.4]
  assign _T_16710 = 7'h2 == _T_10211_63; // @[Mux.scala 46:19:@13525.4]
  assign _T_16711 = _T_16710 ? _T_9260_1 : _T_16709; // @[Mux.scala 46:16:@13526.4]
  assign _T_16712 = 7'h1 == _T_10211_63; // @[Mux.scala 46:19:@13527.4]
  assign _T_16713 = _T_16712 ? _T_9260_0 : _T_16711; // @[Mux.scala 46:16:@13528.4]
  assign _GEN_224 = _T_9256 ? _T_9535_0 : _T_16855_0; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_225 = _T_9256 ? _T_9535_1 : _T_16855_1; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_226 = _T_9256 ? _T_9535_2 : _T_16855_2; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_227 = _T_9256 ? _T_9535_3 : _T_16855_3; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_228 = _T_9256 ? _T_9535_4 : _T_16855_4; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_229 = _T_9256 ? _T_9535_5 : _T_16855_5; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_230 = _T_9256 ? _T_9535_6 : _T_16855_6; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_231 = _T_9256 ? _T_9535_7 : _T_16855_7; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_232 = _T_9256 ? _T_9535_8 : _T_16855_8; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_233 = _T_9256 ? _T_9535_9 : _T_16855_9; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_234 = _T_9256 ? _T_9535_10 : _T_16855_10; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_235 = _T_9256 ? _T_9535_11 : _T_16855_11; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_236 = _T_9256 ? _T_9535_12 : _T_16855_12; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_237 = _T_9256 ? _T_9535_13 : _T_16855_13; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_238 = _T_9256 ? _T_9535_14 : _T_16855_14; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_239 = _T_9256 ? _T_9535_15 : _T_16855_15; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_240 = _T_9256 ? _T_9535_16 : _T_16855_16; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_241 = _T_9256 ? _T_9535_17 : _T_16855_17; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_242 = _T_9256 ? _T_9535_18 : _T_16855_18; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_243 = _T_9256 ? _T_9535_19 : _T_16855_19; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_244 = _T_9256 ? _T_9535_20 : _T_16855_20; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_245 = _T_9256 ? _T_9535_21 : _T_16855_21; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_246 = _T_9256 ? _T_9535_22 : _T_16855_22; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_247 = _T_9256 ? _T_9535_23 : _T_16855_23; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_248 = _T_9256 ? _T_9535_24 : _T_16855_24; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_249 = _T_9256 ? _T_9535_25 : _T_16855_25; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_250 = _T_9256 ? _T_9535_26 : _T_16855_26; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_251 = _T_9256 ? _T_9535_27 : _T_16855_27; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_252 = _T_9256 ? _T_9535_28 : _T_16855_28; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_253 = _T_9256 ? _T_9535_29 : _T_16855_29; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_254 = _T_9256 ? _T_9535_30 : _T_16855_30; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_255 = _T_9256 ? _T_9535_31 : _T_16855_31; // @[NV_NVDLA_CSC_WL_dec.scala 124:19:@13567.4]
  assign _GEN_256 = _T_9330_0 ? _T_10413 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13602.6]
  assign _GEN_258 = _T_9330_1 ? _T_10420 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13610.6]
  assign _GEN_260 = _T_9330_2 ? _T_10430 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13618.6]
  assign _GEN_262 = _T_9330_3 ? _T_10443 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13626.6]
  assign _GEN_264 = _T_9330_4 ? _T_10459 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13634.6]
  assign _GEN_266 = _T_9330_5 ? _T_10478 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13642.6]
  assign _GEN_268 = _T_9330_6 ? _T_10500 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13650.6]
  assign _GEN_270 = _T_9330_7 ? _T_10525 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13658.6]
  assign _GEN_272 = _T_9330_8 ? _T_10553 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13666.6]
  assign _GEN_274 = _T_9330_9 ? _T_10584 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13674.6]
  assign _GEN_276 = _T_9330_10 ? _T_10618 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13682.6]
  assign _GEN_278 = _T_9330_11 ? _T_10655 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13690.6]
  assign _GEN_280 = _T_9330_12 ? _T_10695 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13698.6]
  assign _GEN_282 = _T_9330_13 ? _T_10738 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13706.6]
  assign _GEN_284 = _T_9330_14 ? _T_10784 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13714.6]
  assign _GEN_286 = _T_9330_15 ? _T_10833 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13722.6]
  assign _GEN_288 = _T_9330_16 ? _T_10885 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13730.6]
  assign _GEN_290 = _T_9330_17 ? _T_10940 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13738.6]
  assign _GEN_292 = _T_9330_18 ? _T_10998 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13746.6]
  assign _GEN_294 = _T_9330_19 ? _T_11059 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13754.6]
  assign _GEN_296 = _T_9330_20 ? _T_11123 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13762.6]
  assign _GEN_298 = _T_9330_21 ? _T_11190 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13770.6]
  assign _GEN_300 = _T_9330_22 ? _T_11260 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13778.6]
  assign _GEN_302 = _T_9330_23 ? _T_11333 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13786.6]
  assign _GEN_304 = _T_9330_24 ? _T_11409 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13794.6]
  assign _GEN_306 = _T_9330_25 ? _T_11488 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13802.6]
  assign _GEN_308 = _T_9330_26 ? _T_11570 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13810.6]
  assign _GEN_310 = _T_9330_27 ? _T_11655 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13818.6]
  assign _GEN_312 = _T_9330_28 ? _T_11743 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13826.6]
  assign _GEN_314 = _T_9330_29 ? _T_11834 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13834.6]
  assign _GEN_316 = _T_9330_30 ? _T_11928 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13842.6]
  assign _GEN_318 = _T_9330_31 ? _T_12025 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13850.6]
  assign _GEN_320 = _T_9330_32 ? _T_12125 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13858.6]
  assign _GEN_322 = _T_9330_33 ? _T_12228 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13866.6]
  assign _GEN_324 = _T_9330_34 ? _T_12334 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13874.6]
  assign _GEN_326 = _T_9330_35 ? _T_12443 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13882.6]
  assign _GEN_328 = _T_9330_36 ? _T_12555 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13890.6]
  assign _GEN_330 = _T_9330_37 ? _T_12670 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13898.6]
  assign _GEN_332 = _T_9330_38 ? _T_12788 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13906.6]
  assign _GEN_334 = _T_9330_39 ? _T_12909 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13914.6]
  assign _GEN_336 = _T_9330_40 ? _T_13033 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13922.6]
  assign _GEN_338 = _T_9330_41 ? _T_13160 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13930.6]
  assign _GEN_340 = _T_9330_42 ? _T_13290 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13938.6]
  assign _GEN_342 = _T_9330_43 ? _T_13423 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13946.6]
  assign _GEN_344 = _T_9330_44 ? _T_13559 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13954.6]
  assign _GEN_346 = _T_9330_45 ? _T_13698 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13962.6]
  assign _GEN_348 = _T_9330_46 ? _T_13840 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13970.6]
  assign _GEN_350 = _T_9330_47 ? _T_13985 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13978.6]
  assign _GEN_352 = _T_9330_48 ? _T_14133 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13986.6]
  assign _GEN_354 = _T_9330_49 ? _T_14284 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@13994.6]
  assign _GEN_356 = _T_9330_50 ? _T_14438 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14002.6]
  assign _GEN_358 = _T_9330_51 ? _T_14595 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14010.6]
  assign _GEN_360 = _T_9330_52 ? _T_14755 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14018.6]
  assign _GEN_362 = _T_9330_53 ? _T_14918 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14026.6]
  assign _GEN_364 = _T_9330_54 ? _T_15084 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14034.6]
  assign _GEN_366 = _T_9330_55 ? _T_15253 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14042.6]
  assign _GEN_368 = _T_9330_56 ? _T_15425 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14050.6]
  assign _GEN_370 = _T_9330_57 ? _T_15600 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14058.6]
  assign _GEN_372 = _T_9330_58 ? _T_15778 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14066.6]
  assign _GEN_374 = _T_9330_59 ? _T_15959 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14074.6]
  assign _GEN_376 = _T_9330_60 ? _T_16143 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14082.6]
  assign _GEN_378 = _T_9330_61 ? _T_16330 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14090.6]
  assign _GEN_380 = _T_9330_62 ? _T_16520 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14098.6]
  assign _GEN_382 = _T_9330_63 ? _T_16713 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 129:29:@14106.6]
  assign _T_17161 = _T_10413 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14114.4]
  assign _T_17163 = _T_10420 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14116.4]
  assign _T_17165 = _T_10430 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14118.4]
  assign _T_17167 = _T_10443 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14120.4]
  assign _T_17169 = _T_10459 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14122.4]
  assign _T_17171 = _T_10478 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14124.4]
  assign _T_17173 = _T_10500 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14126.4]
  assign _T_17175 = _T_10525 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14128.4]
  assign _T_17177 = _T_10553 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14130.4]
  assign _T_17179 = _T_10584 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14132.4]
  assign _T_17181 = _T_10618 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14134.4]
  assign _T_17183 = _T_10655 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14136.4]
  assign _T_17185 = _T_10695 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14138.4]
  assign _T_17187 = _T_10738 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14140.4]
  assign _T_17189 = _T_10784 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14142.4]
  assign _T_17191 = _T_10833 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14144.4]
  assign _T_17193 = _T_10885 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14146.4]
  assign _T_17195 = _T_10940 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14148.4]
  assign _T_17197 = _T_10998 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14150.4]
  assign _T_17199 = _T_11059 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14152.4]
  assign _T_17201 = _T_11123 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14154.4]
  assign _T_17203 = _T_11190 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14156.4]
  assign _T_17205 = _T_11260 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14158.4]
  assign _T_17207 = _T_11333 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14160.4]
  assign _T_17209 = _T_11409 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14162.4]
  assign _T_17211 = _T_11488 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14164.4]
  assign _T_17213 = _T_11570 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14166.4]
  assign _T_17215 = _T_11655 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14168.4]
  assign _T_17217 = _T_11743 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14170.4]
  assign _T_17219 = _T_11834 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14172.4]
  assign _T_17221 = _T_11928 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14174.4]
  assign _T_17223 = _T_12025 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14176.4]
  assign _T_17225 = _T_12125 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14178.4]
  assign _T_17227 = _T_12228 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14180.4]
  assign _T_17229 = _T_12334 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14182.4]
  assign _T_17231 = _T_12443 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14184.4]
  assign _T_17233 = _T_12555 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14186.4]
  assign _T_17235 = _T_12670 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14188.4]
  assign _T_17237 = _T_12788 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14190.4]
  assign _T_17239 = _T_12909 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14192.4]
  assign _T_17241 = _T_13033 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14194.4]
  assign _T_17243 = _T_13160 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14196.4]
  assign _T_17245 = _T_13290 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14198.4]
  assign _T_17247 = _T_13423 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14200.4]
  assign _T_17249 = _T_13559 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14202.4]
  assign _T_17251 = _T_13698 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14204.4]
  assign _T_17253 = _T_13840 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14206.4]
  assign _T_17255 = _T_13985 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14208.4]
  assign _T_17257 = _T_14133 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14210.4]
  assign _T_17259 = _T_14284 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14212.4]
  assign _T_17261 = _T_14438 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14214.4]
  assign _T_17263 = _T_14595 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14216.4]
  assign _T_17265 = _T_14755 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14218.4]
  assign _T_17267 = _T_14918 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14220.4]
  assign _T_17269 = _T_15084 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14222.4]
  assign _T_17271 = _T_15253 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14224.4]
  assign _T_17273 = _T_15425 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14226.4]
  assign _T_17275 = _T_15600 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14228.4]
  assign _T_17277 = _T_15778 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14230.4]
  assign _T_17279 = _T_15959 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14232.4]
  assign _T_17281 = _T_16143 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14234.4]
  assign _T_17283 = _T_16330 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14236.4]
  assign _T_17285 = _T_16520 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14238.4]
  assign _T_17287 = _T_16713 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 142:49:@14240.4]
  assign _GEN_448 = _T_16716 ? _T_16855_0 : _T_17499_0; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_449 = _T_16716 ? _T_16855_1 : _T_17499_1; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_450 = _T_16716 ? _T_16855_2 : _T_17499_2; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_451 = _T_16716 ? _T_16855_3 : _T_17499_3; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_452 = _T_16716 ? _T_16855_4 : _T_17499_4; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_453 = _T_16716 ? _T_16855_5 : _T_17499_5; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_454 = _T_16716 ? _T_16855_6 : _T_17499_6; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_455 = _T_16716 ? _T_16855_7 : _T_17499_7; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_456 = _T_16716 ? _T_16855_8 : _T_17499_8; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_457 = _T_16716 ? _T_16855_9 : _T_17499_9; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_458 = _T_16716 ? _T_16855_10 : _T_17499_10; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_459 = _T_16716 ? _T_16855_11 : _T_17499_11; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_460 = _T_16716 ? _T_16855_12 : _T_17499_12; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_461 = _T_16716 ? _T_16855_13 : _T_17499_13; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_462 = _T_16716 ? _T_16855_14 : _T_17499_14; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_463 = _T_16716 ? _T_16855_15 : _T_17499_15; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_464 = _T_16716 ? _T_16855_16 : _T_17499_16; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_465 = _T_16716 ? _T_16855_17 : _T_17499_17; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_466 = _T_16716 ? _T_16855_18 : _T_17499_18; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_467 = _T_16716 ? _T_16855_19 : _T_17499_19; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_468 = _T_16716 ? _T_16855_20 : _T_17499_20; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_469 = _T_16716 ? _T_16855_21 : _T_17499_21; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_470 = _T_16716 ? _T_16855_22 : _T_17499_22; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_471 = _T_16716 ? _T_16855_23 : _T_17499_23; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_472 = _T_16716 ? _T_16855_24 : _T_17499_24; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_473 = _T_16716 ? _T_16855_25 : _T_17499_25; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_474 = _T_16716 ? _T_16855_26 : _T_17499_26; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_475 = _T_16716 ? _T_16855_27 : _T_17499_27; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_476 = _T_16716 ? _T_16855_28 : _T_17499_28; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_477 = _T_16716 ? _T_16855_29 : _T_17499_29; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_478 = _T_16716 ? _T_16855_30 : _T_17499_30; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _GEN_479 = _T_16716 ? _T_16855_31 : _T_17499_31; // @[NV_NVDLA_CSC_WL_dec.scala 153:19:@14280.4]
  assign _T_17676 = {_T_17294_7,_T_17294_6,_T_17294_5,_T_17294_4,_T_17294_3,_T_17294_2,_T_17294_1,_T_17294_0}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14449.4]
  assign _T_17684 = {_T_17294_15,_T_17294_14,_T_17294_13,_T_17294_12,_T_17294_11,_T_17294_10,_T_17294_9,_T_17294_8,_T_17676}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14457.4]
  assign _T_17691 = {_T_17294_23,_T_17294_22,_T_17294_21,_T_17294_20,_T_17294_19,_T_17294_18,_T_17294_17,_T_17294_16}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14464.4]
  assign _T_17700 = {_T_17294_31,_T_17294_30,_T_17294_29,_T_17294_28,_T_17294_27,_T_17294_26,_T_17294_25,_T_17294_24,_T_17691,_T_17684}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14473.4]
  assign _T_17707 = {_T_17294_39,_T_17294_38,_T_17294_37,_T_17294_36,_T_17294_35,_T_17294_34,_T_17294_33,_T_17294_32}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14480.4]
  assign _T_17715 = {_T_17294_47,_T_17294_46,_T_17294_45,_T_17294_44,_T_17294_43,_T_17294_42,_T_17294_41,_T_17294_40,_T_17707}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14488.4]
  assign _T_17722 = {_T_17294_55,_T_17294_54,_T_17294_53,_T_17294_52,_T_17294_51,_T_17294_50,_T_17294_49,_T_17294_48}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14495.4]
  assign _T_17731 = {_T_17294_63,_T_17294_62,_T_17294_61,_T_17294_60,_T_17294_59,_T_17294_58,_T_17294_57,_T_17294_56,_T_17722,_T_17715}; // @[NV_NVDLA_CSC_WL_dec.scala 161:36:@14504.4]
  assign _T_17739 = {_T_17499_7,_T_17499_6,_T_17499_5,_T_17499_4,_T_17499_3,_T_17499_2,_T_17499_1,_T_17499_0}; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14513.4]
  assign _T_17747 = {_T_17499_15,_T_17499_14,_T_17499_13,_T_17499_12,_T_17499_11,_T_17499_10,_T_17499_9,_T_17499_8,_T_17739}; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14521.4]
  assign _T_17754 = {_T_17499_23,_T_17499_22,_T_17499_21,_T_17499_20,_T_17499_19,_T_17499_18,_T_17499_17,_T_17499_16}; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14528.4]
  assign _T_17762 = {_T_17499_31,_T_17499_30,_T_17499_29,_T_17499_28,_T_17499_27,_T_17499_26,_T_17499_25,_T_17499_24,_T_17754}; // @[NV_NVDLA_CSC_WL_dec.scala 162:34:@14536.4]
  assign io_output_valid = _T_17290; // @[NV_NVDLA_CSC_WL_dec.scala 160:21:@14442.4]
  assign io_output_bits_mask = {_T_17731,_T_17700}; // @[NV_NVDLA_CSC_WL_dec.scala 161:25:@14506.4]
  assign io_output_bits_data_0 = _T_17603_0; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14539.4]
  assign io_output_bits_data_1 = _T_17603_1; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14540.4]
  assign io_output_bits_data_2 = _T_17603_2; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14541.4]
  assign io_output_bits_data_3 = _T_17603_3; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14542.4]
  assign io_output_bits_data_4 = _T_17603_4; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14543.4]
  assign io_output_bits_data_5 = _T_17603_5; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14544.4]
  assign io_output_bits_data_6 = _T_17603_6; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14545.4]
  assign io_output_bits_data_7 = _T_17603_7; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14546.4]
  assign io_output_bits_data_8 = _T_17603_8; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14547.4]
  assign io_output_bits_data_9 = _T_17603_9; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14548.4]
  assign io_output_bits_data_10 = _T_17603_10; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14549.4]
  assign io_output_bits_data_11 = _T_17603_11; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14550.4]
  assign io_output_bits_data_12 = _T_17603_12; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14551.4]
  assign io_output_bits_data_13 = _T_17603_13; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14552.4]
  assign io_output_bits_data_14 = _T_17603_14; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14553.4]
  assign io_output_bits_data_15 = _T_17603_15; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14554.4]
  assign io_output_bits_data_16 = _T_17603_16; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14555.4]
  assign io_output_bits_data_17 = _T_17603_17; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14556.4]
  assign io_output_bits_data_18 = _T_17603_18; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14557.4]
  assign io_output_bits_data_19 = _T_17603_19; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14558.4]
  assign io_output_bits_data_20 = _T_17603_20; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14559.4]
  assign io_output_bits_data_21 = _T_17603_21; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14560.4]
  assign io_output_bits_data_22 = _T_17603_22; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14561.4]
  assign io_output_bits_data_23 = _T_17603_23; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14562.4]
  assign io_output_bits_data_24 = _T_17603_24; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14563.4]
  assign io_output_bits_data_25 = _T_17603_25; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14564.4]
  assign io_output_bits_data_26 = _T_17603_26; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14565.4]
  assign io_output_bits_data_27 = _T_17603_27; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14566.4]
  assign io_output_bits_data_28 = _T_17603_28; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14567.4]
  assign io_output_bits_data_29 = _T_17603_29; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14568.4]
  assign io_output_bits_data_30 = _T_17603_30; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14569.4]
  assign io_output_bits_data_31 = _T_17603_31; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14570.4]
  assign io_output_bits_data_32 = _T_17603_32; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14571.4]
  assign io_output_bits_data_33 = _T_17603_33; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14572.4]
  assign io_output_bits_data_34 = _T_17603_34; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14573.4]
  assign io_output_bits_data_35 = _T_17603_35; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14574.4]
  assign io_output_bits_data_36 = _T_17603_36; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14575.4]
  assign io_output_bits_data_37 = _T_17603_37; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14576.4]
  assign io_output_bits_data_38 = _T_17603_38; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14577.4]
  assign io_output_bits_data_39 = _T_17603_39; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14578.4]
  assign io_output_bits_data_40 = _T_17603_40; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14579.4]
  assign io_output_bits_data_41 = _T_17603_41; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14580.4]
  assign io_output_bits_data_42 = _T_17603_42; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14581.4]
  assign io_output_bits_data_43 = _T_17603_43; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14582.4]
  assign io_output_bits_data_44 = _T_17603_44; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14583.4]
  assign io_output_bits_data_45 = _T_17603_45; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14584.4]
  assign io_output_bits_data_46 = _T_17603_46; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14585.4]
  assign io_output_bits_data_47 = _T_17603_47; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14586.4]
  assign io_output_bits_data_48 = _T_17603_48; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14587.4]
  assign io_output_bits_data_49 = _T_17603_49; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14588.4]
  assign io_output_bits_data_50 = _T_17603_50; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14589.4]
  assign io_output_bits_data_51 = _T_17603_51; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14590.4]
  assign io_output_bits_data_52 = _T_17603_52; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14591.4]
  assign io_output_bits_data_53 = _T_17603_53; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14592.4]
  assign io_output_bits_data_54 = _T_17603_54; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14593.4]
  assign io_output_bits_data_55 = _T_17603_55; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14594.4]
  assign io_output_bits_data_56 = _T_17603_56; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14595.4]
  assign io_output_bits_data_57 = _T_17603_57; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14596.4]
  assign io_output_bits_data_58 = _T_17603_58; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14597.4]
  assign io_output_bits_data_59 = _T_17603_59; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14598.4]
  assign io_output_bits_data_60 = _T_17603_60; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14599.4]
  assign io_output_bits_data_61 = _T_17603_61; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14600.4]
  assign io_output_bits_data_62 = _T_17603_62; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14601.4]
  assign io_output_bits_data_63 = _T_17603_63; // @[NV_NVDLA_CSC_WL_dec.scala 163:25:@14602.4]
  assign io_output_bits_sel = {_T_17762,_T_17747}; // @[NV_NVDLA_CSC_WL_dec.scala 162:24:@14538.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_9256 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_9260_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_9260_1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_9260_2 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_9260_3 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_9260_4 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_9260_5 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_9260_6 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_9260_7 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9260_8 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_9260_9 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_9260_10 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_9260_11 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_9260_12 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_9260_13 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_9260_14 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_9260_15 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_9260_16 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_9260_17 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_9260_18 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_9260_19 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_9260_20 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_9260_21 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_9260_22 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_9260_23 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_9260_24 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_9260_25 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_9260_26 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_9260_27 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_9260_28 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_9260_29 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_9260_30 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_9260_31 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_9260_32 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_9260_33 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_9260_34 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_9260_35 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_9260_36 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_9260_37 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_9260_38 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_9260_39 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_9260_40 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_9260_41 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_9260_42 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_9260_43 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_9260_44 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_9260_45 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_9260_46 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_9260_47 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_9260_48 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_9260_49 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_9260_50 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_9260_51 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_9260_52 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_9260_53 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_9260_54 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_9260_55 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_9260_56 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_9260_57 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_9260_58 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_9260_59 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_9260_60 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_9260_61 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_9260_62 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_9260_63 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_9330_0 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_9330_1 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_9330_2 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_9330_3 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_9330_4 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_9330_5 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_9330_6 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_9330_7 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_9330_8 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_9330_9 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_9330_10 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_9330_11 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_9330_12 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_9330_13 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_9330_14 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_9330_15 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_9330_16 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_9330_17 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_9330_18 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_9330_19 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_9330_20 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_9330_21 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_9330_22 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_9330_23 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_9330_24 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_9330_25 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_9330_26 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_9330_27 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_9330_28 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_9330_29 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_9330_30 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_9330_31 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_9330_32 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_9330_33 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_9330_34 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_9330_35 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_9330_36 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_9330_37 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_9330_38 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_9330_39 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_9330_40 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_9330_41 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_9330_42 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_9330_43 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_9330_44 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_9330_45 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_9330_46 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_9330_47 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_9330_48 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_9330_49 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_9330_50 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_9330_51 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_9330_52 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_9330_53 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_9330_54 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_9330_55 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_9330_56 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_9330_57 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_9330_58 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_9330_59 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_9330_60 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_9330_61 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_9330_62 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_9330_63 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_9535_0 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_9535_1 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_9535_2 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_9535_3 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_9535_4 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_9535_5 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_9535_6 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_9535_7 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_9535_8 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_9535_9 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_9535_10 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_9535_11 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_9535_12 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_9535_13 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_9535_14 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_9535_15 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_9535_16 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_9535_17 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_9535_18 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_9535_19 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_9535_20 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_9535_21 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_9535_22 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_9535_23 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_9535_24 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_9535_25 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_9535_26 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_9535_27 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_9535_28 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_9535_29 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_9535_30 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_9535_31 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_10211_63 = _RAND_161[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_10211_62 = _RAND_162[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_10211_61 = _RAND_163[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_10211_60 = _RAND_164[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_10211_59 = _RAND_165[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_10211_58 = _RAND_166[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_10211_57 = _RAND_167[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_10211_56 = _RAND_168[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_10211_55 = _RAND_169[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_10211_54 = _RAND_170[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_10211_53 = _RAND_171[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_10211_52 = _RAND_172[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_10211_51 = _RAND_173[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_10211_50 = _RAND_174[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_10211_49 = _RAND_175[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_10211_48 = _RAND_176[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_10211_47 = _RAND_177[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_10211_46 = _RAND_178[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_10211_45 = _RAND_179[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_10211_44 = _RAND_180[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_10211_43 = _RAND_181[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_10211_42 = _RAND_182[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_10211_41 = _RAND_183[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_10211_40 = _RAND_184[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_10211_39 = _RAND_185[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_10211_38 = _RAND_186[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_10211_37 = _RAND_187[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_10211_36 = _RAND_188[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_10211_35 = _RAND_189[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_10211_34 = _RAND_190[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_10211_33 = _RAND_191[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_10211_32 = _RAND_192[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_10211_31 = _RAND_193[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_10211_30 = _RAND_194[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_10211_29 = _RAND_195[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_10211_28 = _RAND_196[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_10211_27 = _RAND_197[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_10211_26 = _RAND_198[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_10211_25 = _RAND_199[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_10211_24 = _RAND_200[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_10211_23 = _RAND_201[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_10211_22 = _RAND_202[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_10211_21 = _RAND_203[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_10211_20 = _RAND_204[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_10211_19 = _RAND_205[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_10211_18 = _RAND_206[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_10211_17 = _RAND_207[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_10211_16 = _RAND_208[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_10211_15 = _RAND_209[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_10211_14 = _RAND_210[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_10211_13 = _RAND_211[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_10211_12 = _RAND_212[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_10211_11 = _RAND_213[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_10211_10 = _RAND_214[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_10211_9 = _RAND_215[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_10211_8 = _RAND_216[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_10211_7 = _RAND_217[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_10211_6 = _RAND_218[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_10211_5 = _RAND_219[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_10211_4 = _RAND_220[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_10211_3 = _RAND_221[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_10211_2 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_10211_1 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_10211_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_16716 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_16855_0 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_16855_1 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_16855_2 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_16855_3 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_16855_4 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_16855_5 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_16855_6 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_16855_7 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_16855_8 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_16855_9 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_16855_10 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_16855_11 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_16855_12 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_16855_13 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_16855_14 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_16855_15 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_16855_16 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_16855_17 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_16855_18 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_16855_19 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_16855_20 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_16855_21 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_16855_22 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_16855_23 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_16855_24 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_16855_25 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_16855_26 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_16855_27 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_16855_28 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_16855_29 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_16855_30 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_16855_31 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_16959_0 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_16959_1 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_16959_2 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_16959_3 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_16959_4 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_16959_5 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_16959_6 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_16959_7 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_16959_8 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_16959_9 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_16959_10 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_16959_11 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_16959_12 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_16959_13 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_16959_14 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_16959_15 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_16959_16 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_16959_17 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_16959_18 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_16959_19 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_16959_20 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_16959_21 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_16959_22 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_16959_23 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_16959_24 = _RAND_282[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_16959_25 = _RAND_283[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_16959_26 = _RAND_284[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_16959_27 = _RAND_285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_16959_28 = _RAND_286[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_16959_29 = _RAND_287[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_16959_30 = _RAND_288[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_16959_31 = _RAND_289[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_16959_32 = _RAND_290[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_16959_33 = _RAND_291[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_16959_34 = _RAND_292[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_16959_35 = _RAND_293[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_16959_36 = _RAND_294[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_16959_37 = _RAND_295[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_16959_38 = _RAND_296[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_16959_39 = _RAND_297[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_16959_40 = _RAND_298[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_16959_41 = _RAND_299[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_16959_42 = _RAND_300[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_16959_43 = _RAND_301[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_16959_44 = _RAND_302[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_16959_45 = _RAND_303[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_16959_46 = _RAND_304[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_16959_47 = _RAND_305[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_16959_48 = _RAND_306[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_16959_49 = _RAND_307[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_16959_50 = _RAND_308[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_16959_51 = _RAND_309[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_16959_52 = _RAND_310[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_16959_53 = _RAND_311[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_16959_54 = _RAND_312[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_16959_55 = _RAND_313[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_16959_56 = _RAND_314[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_16959_57 = _RAND_315[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_16959_58 = _RAND_316[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_16959_59 = _RAND_317[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_16959_60 = _RAND_318[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_16959_61 = _RAND_319[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_16959_62 = _RAND_320[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_16959_63 = _RAND_321[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_17290 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_17294_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_17294_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_17294_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_17294_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_17294_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_17294_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_17294_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_17294_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_17294_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_17294_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_17294_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_17294_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_17294_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_17294_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_17294_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_17294_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_17294_16 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_17294_17 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_17294_18 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_17294_19 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_17294_20 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_17294_21 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_17294_22 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_17294_23 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_17294_24 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_17294_25 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_17294_26 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_17294_27 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_17294_28 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_17294_29 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_17294_30 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_17294_31 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_17294_32 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_17294_33 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_17294_34 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_17294_35 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_17294_36 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_17294_37 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_17294_38 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_17294_39 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_17294_40 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_17294_41 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_17294_42 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_17294_43 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_17294_44 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_17294_45 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_17294_46 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_17294_47 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_17294_48 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_17294_49 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_17294_50 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_17294_51 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_17294_52 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_17294_53 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_17294_54 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_17294_55 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_17294_56 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_17294_57 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_17294_58 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_17294_59 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_17294_60 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_17294_61 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_17294_62 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_17294_63 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_17499_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_17499_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_17499_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_17499_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_17499_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_17499_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_17499_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_17499_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_17499_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_17499_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_17499_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_17499_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_17499_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_17499_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_17499_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_17499_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_17499_16 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_17499_17 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_17499_18 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_17499_19 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_17499_20 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_17499_21 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_17499_22 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_17499_23 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_17499_24 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_17499_25 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_17499_26 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_17499_27 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_17499_28 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_17499_29 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_17499_30 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_17499_31 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_17603_0 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_17603_1 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_17603_2 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_17603_3 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_17603_4 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_17603_5 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_17603_6 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_17603_7 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_17603_8 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_17603_9 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_17603_10 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_17603_11 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_17603_12 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_17603_13 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_17603_14 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_17603_15 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_17603_16 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_17603_17 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_17603_18 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_17603_19 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_17603_20 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_17603_21 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_17603_22 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_17603_23 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_17603_24 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_17603_25 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_17603_26 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_17603_27 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_17603_28 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_17603_29 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_17603_30 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_17603_31 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_17603_32 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_17603_33 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_17603_34 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_17603_35 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_17603_36 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_17603_37 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_17603_38 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_17603_39 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_17603_40 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_17603_41 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_17603_42 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_17603_43 = _RAND_462[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_17603_44 = _RAND_463[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_17603_45 = _RAND_464[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_17603_46 = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_17603_47 = _RAND_466[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_17603_48 = _RAND_467[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_17603_49 = _RAND_468[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_17603_50 = _RAND_469[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_17603_51 = _RAND_470[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_17603_52 = _RAND_471[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_17603_53 = _RAND_472[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_17603_54 = _RAND_473[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_17603_55 = _RAND_474[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_17603_56 = _RAND_475[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_17603_57 = _RAND_476[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_17603_58 = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_17603_59 = _RAND_478[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_17603_60 = _RAND_479[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_17603_61 = _RAND_480[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_17603_62 = _RAND_481[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_17603_63 = _RAND_482[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (_T_326) begin
      _T_9256 <= 1'h0;
    end else begin
      _T_9256 <= io_input_valid;
    end
    if (io_input_valid) begin
      _T_9260_0 <= _T_531;
    end
    if (io_input_valid) begin
      _T_9260_1 <= _T_532;
    end
    if (io_input_valid) begin
      _T_9260_2 <= _T_533;
    end
    if (io_input_valid) begin
      _T_9260_3 <= _T_534;
    end
    if (io_input_valid) begin
      _T_9260_4 <= _T_535;
    end
    if (io_input_valid) begin
      _T_9260_5 <= _T_536;
    end
    if (io_input_valid) begin
      _T_9260_6 <= _T_537;
    end
    if (io_input_valid) begin
      _T_9260_7 <= _T_538;
    end
    if (io_input_valid) begin
      _T_9260_8 <= _T_539;
    end
    if (io_input_valid) begin
      _T_9260_9 <= _T_540;
    end
    if (io_input_valid) begin
      _T_9260_10 <= _T_541;
    end
    if (io_input_valid) begin
      _T_9260_11 <= _T_542;
    end
    if (io_input_valid) begin
      _T_9260_12 <= _T_543;
    end
    if (io_input_valid) begin
      _T_9260_13 <= _T_544;
    end
    if (io_input_valid) begin
      _T_9260_14 <= _T_545;
    end
    if (io_input_valid) begin
      _T_9260_15 <= _T_546;
    end
    if (io_input_valid) begin
      _T_9260_16 <= _T_547;
    end
    if (io_input_valid) begin
      _T_9260_17 <= _T_548;
    end
    if (io_input_valid) begin
      _T_9260_18 <= _T_549;
    end
    if (io_input_valid) begin
      _T_9260_19 <= _T_550;
    end
    if (io_input_valid) begin
      _T_9260_20 <= _T_551;
    end
    if (io_input_valid) begin
      _T_9260_21 <= _T_552;
    end
    if (io_input_valid) begin
      _T_9260_22 <= _T_553;
    end
    if (io_input_valid) begin
      _T_9260_23 <= _T_554;
    end
    if (io_input_valid) begin
      _T_9260_24 <= _T_555;
    end
    if (io_input_valid) begin
      _T_9260_25 <= _T_556;
    end
    if (io_input_valid) begin
      _T_9260_26 <= _T_557;
    end
    if (io_input_valid) begin
      _T_9260_27 <= _T_558;
    end
    if (io_input_valid) begin
      _T_9260_28 <= _T_559;
    end
    if (io_input_valid) begin
      _T_9260_29 <= _T_560;
    end
    if (io_input_valid) begin
      _T_9260_30 <= _T_561;
    end
    if (io_input_valid) begin
      _T_9260_31 <= _T_562;
    end
    if (io_input_valid) begin
      _T_9260_32 <= _T_563;
    end
    if (io_input_valid) begin
      _T_9260_33 <= _T_564;
    end
    if (io_input_valid) begin
      _T_9260_34 <= _T_565;
    end
    if (io_input_valid) begin
      _T_9260_35 <= _T_566;
    end
    if (io_input_valid) begin
      _T_9260_36 <= _T_567;
    end
    if (io_input_valid) begin
      _T_9260_37 <= _T_568;
    end
    if (io_input_valid) begin
      _T_9260_38 <= _T_569;
    end
    if (io_input_valid) begin
      _T_9260_39 <= _T_570;
    end
    if (io_input_valid) begin
      _T_9260_40 <= _T_571;
    end
    if (io_input_valid) begin
      _T_9260_41 <= _T_572;
    end
    if (io_input_valid) begin
      _T_9260_42 <= _T_573;
    end
    if (io_input_valid) begin
      _T_9260_43 <= _T_574;
    end
    if (io_input_valid) begin
      _T_9260_44 <= _T_575;
    end
    if (io_input_valid) begin
      _T_9260_45 <= _T_576;
    end
    if (io_input_valid) begin
      _T_9260_46 <= _T_577;
    end
    if (io_input_valid) begin
      _T_9260_47 <= _T_578;
    end
    if (io_input_valid) begin
      _T_9260_48 <= _T_579;
    end
    if (io_input_valid) begin
      _T_9260_49 <= _T_580;
    end
    if (io_input_valid) begin
      _T_9260_50 <= _T_581;
    end
    if (io_input_valid) begin
      _T_9260_51 <= _T_582;
    end
    if (io_input_valid) begin
      _T_9260_52 <= _T_583;
    end
    if (io_input_valid) begin
      _T_9260_53 <= _T_584;
    end
    if (io_input_valid) begin
      _T_9260_54 <= _T_585;
    end
    if (io_input_valid) begin
      _T_9260_55 <= _T_586;
    end
    if (io_input_valid) begin
      _T_9260_56 <= _T_587;
    end
    if (io_input_valid) begin
      _T_9260_57 <= _T_588;
    end
    if (io_input_valid) begin
      _T_9260_58 <= _T_589;
    end
    if (io_input_valid) begin
      _T_9260_59 <= _T_590;
    end
    if (io_input_valid) begin
      _T_9260_60 <= _T_591;
    end
    if (io_input_valid) begin
      _T_9260_61 <= _T_592;
    end
    if (io_input_valid) begin
      _T_9260_62 <= _T_593;
    end
    if (io_input_valid) begin
      _T_9260_63 <= _T_594;
    end
    if (io_input_valid) begin
      _T_9330_0 <= _T_397;
    end
    if (io_input_valid) begin
      _T_9330_1 <= _T_398;
    end
    if (io_input_valid) begin
      _T_9330_2 <= _T_399;
    end
    if (io_input_valid) begin
      _T_9330_3 <= _T_400;
    end
    if (io_input_valid) begin
      _T_9330_4 <= _T_401;
    end
    if (io_input_valid) begin
      _T_9330_5 <= _T_402;
    end
    if (io_input_valid) begin
      _T_9330_6 <= _T_403;
    end
    if (io_input_valid) begin
      _T_9330_7 <= _T_404;
    end
    if (io_input_valid) begin
      _T_9330_8 <= _T_405;
    end
    if (io_input_valid) begin
      _T_9330_9 <= _T_406;
    end
    if (io_input_valid) begin
      _T_9330_10 <= _T_407;
    end
    if (io_input_valid) begin
      _T_9330_11 <= _T_408;
    end
    if (io_input_valid) begin
      _T_9330_12 <= _T_409;
    end
    if (io_input_valid) begin
      _T_9330_13 <= _T_410;
    end
    if (io_input_valid) begin
      _T_9330_14 <= _T_411;
    end
    if (io_input_valid) begin
      _T_9330_15 <= _T_412;
    end
    if (io_input_valid) begin
      _T_9330_16 <= _T_413;
    end
    if (io_input_valid) begin
      _T_9330_17 <= _T_414;
    end
    if (io_input_valid) begin
      _T_9330_18 <= _T_415;
    end
    if (io_input_valid) begin
      _T_9330_19 <= _T_416;
    end
    if (io_input_valid) begin
      _T_9330_20 <= _T_417;
    end
    if (io_input_valid) begin
      _T_9330_21 <= _T_418;
    end
    if (io_input_valid) begin
      _T_9330_22 <= _T_419;
    end
    if (io_input_valid) begin
      _T_9330_23 <= _T_420;
    end
    if (io_input_valid) begin
      _T_9330_24 <= _T_421;
    end
    if (io_input_valid) begin
      _T_9330_25 <= _T_422;
    end
    if (io_input_valid) begin
      _T_9330_26 <= _T_423;
    end
    if (io_input_valid) begin
      _T_9330_27 <= _T_424;
    end
    if (io_input_valid) begin
      _T_9330_28 <= _T_425;
    end
    if (io_input_valid) begin
      _T_9330_29 <= _T_426;
    end
    if (io_input_valid) begin
      _T_9330_30 <= _T_427;
    end
    if (io_input_valid) begin
      _T_9330_31 <= _T_428;
    end
    if (io_input_valid) begin
      _T_9330_32 <= _T_429;
    end
    if (io_input_valid) begin
      _T_9330_33 <= _T_430;
    end
    if (io_input_valid) begin
      _T_9330_34 <= _T_431;
    end
    if (io_input_valid) begin
      _T_9330_35 <= _T_432;
    end
    if (io_input_valid) begin
      _T_9330_36 <= _T_433;
    end
    if (io_input_valid) begin
      _T_9330_37 <= _T_434;
    end
    if (io_input_valid) begin
      _T_9330_38 <= _T_435;
    end
    if (io_input_valid) begin
      _T_9330_39 <= _T_436;
    end
    if (io_input_valid) begin
      _T_9330_40 <= _T_437;
    end
    if (io_input_valid) begin
      _T_9330_41 <= _T_438;
    end
    if (io_input_valid) begin
      _T_9330_42 <= _T_439;
    end
    if (io_input_valid) begin
      _T_9330_43 <= _T_440;
    end
    if (io_input_valid) begin
      _T_9330_44 <= _T_441;
    end
    if (io_input_valid) begin
      _T_9330_45 <= _T_442;
    end
    if (io_input_valid) begin
      _T_9330_46 <= _T_443;
    end
    if (io_input_valid) begin
      _T_9330_47 <= _T_444;
    end
    if (io_input_valid) begin
      _T_9330_48 <= _T_445;
    end
    if (io_input_valid) begin
      _T_9330_49 <= _T_446;
    end
    if (io_input_valid) begin
      _T_9330_50 <= _T_447;
    end
    if (io_input_valid) begin
      _T_9330_51 <= _T_448;
    end
    if (io_input_valid) begin
      _T_9330_52 <= _T_449;
    end
    if (io_input_valid) begin
      _T_9330_53 <= _T_450;
    end
    if (io_input_valid) begin
      _T_9330_54 <= _T_451;
    end
    if (io_input_valid) begin
      _T_9330_55 <= _T_452;
    end
    if (io_input_valid) begin
      _T_9330_56 <= _T_453;
    end
    if (io_input_valid) begin
      _T_9330_57 <= _T_454;
    end
    if (io_input_valid) begin
      _T_9330_58 <= _T_455;
    end
    if (io_input_valid) begin
      _T_9330_59 <= _T_456;
    end
    if (io_input_valid) begin
      _T_9330_60 <= _T_457;
    end
    if (io_input_valid) begin
      _T_9330_61 <= _T_458;
    end
    if (io_input_valid) begin
      _T_9330_62 <= _T_459;
    end
    if (io_input_valid) begin
      _T_9330_63 <= _T_460;
    end
    if (_T_326) begin
      _T_9535_0 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_0 <= _T_633;
      end
    end
    if (_T_326) begin
      _T_9535_1 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_1 <= _T_634;
      end
    end
    if (_T_326) begin
      _T_9535_2 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_2 <= _T_635;
      end
    end
    if (_T_326) begin
      _T_9535_3 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_3 <= _T_636;
      end
    end
    if (_T_326) begin
      _T_9535_4 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_4 <= _T_637;
      end
    end
    if (_T_326) begin
      _T_9535_5 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_5 <= _T_638;
      end
    end
    if (_T_326) begin
      _T_9535_6 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_6 <= _T_639;
      end
    end
    if (_T_326) begin
      _T_9535_7 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_7 <= _T_640;
      end
    end
    if (_T_326) begin
      _T_9535_8 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_8 <= _T_641;
      end
    end
    if (_T_326) begin
      _T_9535_9 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_9 <= _T_642;
      end
    end
    if (_T_326) begin
      _T_9535_10 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_10 <= _T_643;
      end
    end
    if (_T_326) begin
      _T_9535_11 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_11 <= _T_644;
      end
    end
    if (_T_326) begin
      _T_9535_12 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_12 <= _T_645;
      end
    end
    if (_T_326) begin
      _T_9535_13 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_13 <= _T_646;
      end
    end
    if (_T_326) begin
      _T_9535_14 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_14 <= _T_647;
      end
    end
    if (_T_326) begin
      _T_9535_15 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_15 <= _T_648;
      end
    end
    if (_T_326) begin
      _T_9535_16 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_16 <= _T_649;
      end
    end
    if (_T_326) begin
      _T_9535_17 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_17 <= _T_650;
      end
    end
    if (_T_326) begin
      _T_9535_18 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_18 <= _T_651;
      end
    end
    if (_T_326) begin
      _T_9535_19 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_19 <= _T_652;
      end
    end
    if (_T_326) begin
      _T_9535_20 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_20 <= _T_653;
      end
    end
    if (_T_326) begin
      _T_9535_21 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_21 <= _T_654;
      end
    end
    if (_T_326) begin
      _T_9535_22 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_22 <= _T_655;
      end
    end
    if (_T_326) begin
      _T_9535_23 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_23 <= _T_656;
      end
    end
    if (_T_326) begin
      _T_9535_24 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_24 <= _T_657;
      end
    end
    if (_T_326) begin
      _T_9535_25 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_25 <= _T_658;
      end
    end
    if (_T_326) begin
      _T_9535_26 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_26 <= _T_659;
      end
    end
    if (_T_326) begin
      _T_9535_27 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_27 <= _T_660;
      end
    end
    if (_T_326) begin
      _T_9535_28 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_28 <= _T_661;
      end
    end
    if (_T_326) begin
      _T_9535_29 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_29 <= _T_662;
      end
    end
    if (_T_326) begin
      _T_9535_30 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_30 <= _T_663;
      end
    end
    if (_T_326) begin
      _T_9535_31 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_9535_31 <= _T_664;
      end
    end
    if (_T_326) begin
      _T_10211_63 <= 7'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_63 <= _T_9253;
      end
    end
    if (_T_326) begin
      _T_10211_62 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_62 <= _T_1061_62;
      end
    end
    if (_T_326) begin
      _T_10211_61 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_61 <= _T_1061_61;
      end
    end
    if (_T_326) begin
      _T_10211_60 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_60 <= _T_1061_60;
      end
    end
    if (_T_326) begin
      _T_10211_59 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_59 <= _T_1061_59;
      end
    end
    if (_T_326) begin
      _T_10211_58 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_58 <= _T_1061_58;
      end
    end
    if (_T_326) begin
      _T_10211_57 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_57 <= _T_1061_57;
      end
    end
    if (_T_326) begin
      _T_10211_56 <= 6'h0;
    end else begin
      if (_T_10325) begin
        _T_10211_56 <= _T_1061_56;
      end
    end
    if (_T_326) begin
      _T_10211_55 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_55 <= _T_1061_55;
      end
    end
    if (_T_326) begin
      _T_10211_54 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_54 <= _T_1061_54;
      end
    end
    if (_T_326) begin
      _T_10211_53 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_53 <= _T_1061_53;
      end
    end
    if (_T_326) begin
      _T_10211_52 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_52 <= _T_1061_52;
      end
    end
    if (_T_326) begin
      _T_10211_51 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_51 <= _T_1061_51;
      end
    end
    if (_T_326) begin
      _T_10211_50 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_50 <= _T_1061_50;
      end
    end
    if (_T_326) begin
      _T_10211_49 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_49 <= _T_1061_49;
      end
    end
    if (_T_326) begin
      _T_10211_48 <= 6'h0;
    end else begin
      if (_T_10309) begin
        _T_10211_48 <= _T_1061_48;
      end
    end
    if (_T_326) begin
      _T_10211_47 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_47 <= _T_1061_47;
      end
    end
    if (_T_326) begin
      _T_10211_46 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_46 <= _T_1061_46;
      end
    end
    if (_T_326) begin
      _T_10211_45 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_45 <= _T_1061_45;
      end
    end
    if (_T_326) begin
      _T_10211_44 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_44 <= _T_1061_44;
      end
    end
    if (_T_326) begin
      _T_10211_43 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_43 <= _T_1061_43;
      end
    end
    if (_T_326) begin
      _T_10211_42 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_42 <= _T_1061_42;
      end
    end
    if (_T_326) begin
      _T_10211_41 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_41 <= _T_1061_41;
      end
    end
    if (_T_326) begin
      _T_10211_40 <= 6'h0;
    end else begin
      if (_T_10293) begin
        _T_10211_40 <= _T_1061_40;
      end
    end
    if (_T_326) begin
      _T_10211_39 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_39 <= _T_1061_39;
      end
    end
    if (_T_326) begin
      _T_10211_38 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_38 <= _T_1061_38;
      end
    end
    if (_T_326) begin
      _T_10211_37 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_37 <= _T_1061_37;
      end
    end
    if (_T_326) begin
      _T_10211_36 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_36 <= _T_1061_36;
      end
    end
    if (_T_326) begin
      _T_10211_35 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_35 <= _T_1061_35;
      end
    end
    if (_T_326) begin
      _T_10211_34 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_34 <= _T_1061_34;
      end
    end
    if (_T_326) begin
      _T_10211_33 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_33 <= _T_1061_33;
      end
    end
    if (_T_326) begin
      _T_10211_32 <= 6'h0;
    end else begin
      if (_T_10277) begin
        _T_10211_32 <= _T_1061_32;
      end
    end
    if (_T_326) begin
      _T_10211_31 <= 6'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_31 <= _T_4133;
      end
    end
    if (_T_326) begin
      _T_10211_30 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_30 <= _T_1061_30;
      end
    end
    if (_T_326) begin
      _T_10211_29 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_29 <= _T_1061_29;
      end
    end
    if (_T_326) begin
      _T_10211_28 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_28 <= _T_1061_28;
      end
    end
    if (_T_326) begin
      _T_10211_27 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_27 <= _T_1061_27;
      end
    end
    if (_T_326) begin
      _T_10211_26 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_26 <= _T_1061_26;
      end
    end
    if (_T_326) begin
      _T_10211_25 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_25 <= _T_1061_25;
      end
    end
    if (_T_326) begin
      _T_10211_24 <= 5'h0;
    end else begin
      if (_T_10261) begin
        _T_10211_24 <= _T_1061_24;
      end
    end
    if (_T_326) begin
      _T_10211_23 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_23 <= _T_1061_23;
      end
    end
    if (_T_326) begin
      _T_10211_22 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_22 <= _T_1061_22;
      end
    end
    if (_T_326) begin
      _T_10211_21 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_21 <= _T_1061_21;
      end
    end
    if (_T_326) begin
      _T_10211_20 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_20 <= _T_1061_20;
      end
    end
    if (_T_326) begin
      _T_10211_19 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_19 <= _T_1061_19;
      end
    end
    if (_T_326) begin
      _T_10211_18 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_18 <= _T_1061_18;
      end
    end
    if (_T_326) begin
      _T_10211_17 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_17 <= _T_1061_17;
      end
    end
    if (_T_326) begin
      _T_10211_16 <= 5'h0;
    end else begin
      if (_T_10245) begin
        _T_10211_16 <= _T_1061_16;
      end
    end
    if (_T_326) begin
      _T_10211_15 <= 5'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_15 <= _T_2341;
      end
    end
    if (_T_326) begin
      _T_10211_14 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_14 <= _T_1061_14;
      end
    end
    if (_T_326) begin
      _T_10211_13 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_13 <= _T_1061_13;
      end
    end
    if (_T_326) begin
      _T_10211_12 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_12 <= _T_1061_12;
      end
    end
    if (_T_326) begin
      _T_10211_11 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_11 <= _T_1061_11;
      end
    end
    if (_T_326) begin
      _T_10211_10 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_10 <= _T_1061_10;
      end
    end
    if (_T_326) begin
      _T_10211_9 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_9 <= _T_1061_9;
      end
    end
    if (_T_326) begin
      _T_10211_8 <= 4'h0;
    end else begin
      if (_T_10229) begin
        _T_10211_8 <= _T_1061_8;
      end
    end
    if (_T_326) begin
      _T_10211_7 <= 4'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_7 <= _T_1637;
      end
    end
    if (_T_326) begin
      _T_10211_6 <= 3'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_6 <= _T_1061_6;
      end
    end
    if (_T_326) begin
      _T_10211_5 <= 3'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_5 <= _T_1061_5;
      end
    end
    if (_T_326) begin
      _T_10211_4 <= 3'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_4 <= _T_1061_4;
      end
    end
    if (_T_326) begin
      _T_10211_3 <= 3'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_3 <= _T_1333;
      end
    end
    if (_T_326) begin
      _T_10211_2 <= 2'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_2 <= _T_1061_2;
      end
    end
    if (_T_326) begin
      _T_10211_1 <= 2'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_1 <= _T_1193;
      end
    end
    if (_T_326) begin
      _T_10211_0 <= 1'h0;
    end else begin
      if (_T_10213) begin
        _T_10211_0 <= _T_1125;
      end
    end
    if (_T_326) begin
      _T_16716 <= 1'h0;
    end else begin
      _T_16716 <= _T_9256;
    end
    if (_T_326) begin
      _T_16855_0 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_0 <= _T_9535_0;
      end
    end
    if (_T_326) begin
      _T_16855_1 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_1 <= _T_9535_1;
      end
    end
    if (_T_326) begin
      _T_16855_2 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_2 <= _T_9535_2;
      end
    end
    if (_T_326) begin
      _T_16855_3 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_3 <= _T_9535_3;
      end
    end
    if (_T_326) begin
      _T_16855_4 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_4 <= _T_9535_4;
      end
    end
    if (_T_326) begin
      _T_16855_5 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_5 <= _T_9535_5;
      end
    end
    if (_T_326) begin
      _T_16855_6 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_6 <= _T_9535_6;
      end
    end
    if (_T_326) begin
      _T_16855_7 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_7 <= _T_9535_7;
      end
    end
    if (_T_326) begin
      _T_16855_8 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_8 <= _T_9535_8;
      end
    end
    if (_T_326) begin
      _T_16855_9 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_9 <= _T_9535_9;
      end
    end
    if (_T_326) begin
      _T_16855_10 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_10 <= _T_9535_10;
      end
    end
    if (_T_326) begin
      _T_16855_11 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_11 <= _T_9535_11;
      end
    end
    if (_T_326) begin
      _T_16855_12 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_12 <= _T_9535_12;
      end
    end
    if (_T_326) begin
      _T_16855_13 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_13 <= _T_9535_13;
      end
    end
    if (_T_326) begin
      _T_16855_14 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_14 <= _T_9535_14;
      end
    end
    if (_T_326) begin
      _T_16855_15 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_15 <= _T_9535_15;
      end
    end
    if (_T_326) begin
      _T_16855_16 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_16 <= _T_9535_16;
      end
    end
    if (_T_326) begin
      _T_16855_17 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_17 <= _T_9535_17;
      end
    end
    if (_T_326) begin
      _T_16855_18 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_18 <= _T_9535_18;
      end
    end
    if (_T_326) begin
      _T_16855_19 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_19 <= _T_9535_19;
      end
    end
    if (_T_326) begin
      _T_16855_20 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_20 <= _T_9535_20;
      end
    end
    if (_T_326) begin
      _T_16855_21 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_21 <= _T_9535_21;
      end
    end
    if (_T_326) begin
      _T_16855_22 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_22 <= _T_9535_22;
      end
    end
    if (_T_326) begin
      _T_16855_23 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_23 <= _T_9535_23;
      end
    end
    if (_T_326) begin
      _T_16855_24 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_24 <= _T_9535_24;
      end
    end
    if (_T_326) begin
      _T_16855_25 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_25 <= _T_9535_25;
      end
    end
    if (_T_326) begin
      _T_16855_26 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_26 <= _T_9535_26;
      end
    end
    if (_T_326) begin
      _T_16855_27 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_27 <= _T_9535_27;
      end
    end
    if (_T_326) begin
      _T_16855_28 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_28 <= _T_9535_28;
      end
    end
    if (_T_326) begin
      _T_16855_29 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_29 <= _T_9535_29;
      end
    end
    if (_T_326) begin
      _T_16855_30 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_30 <= _T_9535_30;
      end
    end
    if (_T_326) begin
      _T_16855_31 <= 1'h0;
    end else begin
      if (_T_9256) begin
        _T_16855_31 <= _T_9535_31;
      end
    end
    if (_T_9256) begin
      if (_T_9330_0) begin
        if (_T_10211_0) begin
          _T_16959_0 <= _T_9260_0;
        end else begin
          _T_16959_0 <= 8'h0;
        end
      end else begin
        _T_16959_0 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_1) begin
        if (_T_10419) begin
          _T_16959_1 <= _T_9260_0;
        end else begin
          if (_T_10417) begin
            _T_16959_1 <= _T_9260_1;
          end else begin
            _T_16959_1 <= 8'h0;
          end
        end
      end else begin
        _T_16959_1 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_2) begin
        if (_T_10429) begin
          _T_16959_2 <= _T_9260_0;
        end else begin
          if (_T_10427) begin
            _T_16959_2 <= _T_9260_1;
          end else begin
            if (_T_10425) begin
              _T_16959_2 <= _T_9260_2;
            end else begin
              _T_16959_2 <= 8'h0;
            end
          end
        end
      end else begin
        _T_16959_2 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_3) begin
        if (_T_10442) begin
          _T_16959_3 <= _T_9260_0;
        end else begin
          if (_T_10440) begin
            _T_16959_3 <= _T_9260_1;
          end else begin
            if (_T_10438) begin
              _T_16959_3 <= _T_9260_2;
            end else begin
              if (_T_10436) begin
                _T_16959_3 <= _T_9260_3;
              end else begin
                _T_16959_3 <= 8'h0;
              end
            end
          end
        end
      end else begin
        _T_16959_3 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_4) begin
        if (_T_10458) begin
          _T_16959_4 <= _T_9260_0;
        end else begin
          if (_T_10456) begin
            _T_16959_4 <= _T_9260_1;
          end else begin
            if (_T_10454) begin
              _T_16959_4 <= _T_9260_2;
            end else begin
              if (_T_10452) begin
                _T_16959_4 <= _T_9260_3;
              end else begin
                if (_T_10450) begin
                  _T_16959_4 <= _T_9260_4;
                end else begin
                  _T_16959_4 <= 8'h0;
                end
              end
            end
          end
        end
      end else begin
        _T_16959_4 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_5) begin
        if (_T_10477) begin
          _T_16959_5 <= _T_9260_0;
        end else begin
          if (_T_10475) begin
            _T_16959_5 <= _T_9260_1;
          end else begin
            if (_T_10473) begin
              _T_16959_5 <= _T_9260_2;
            end else begin
              if (_T_10471) begin
                _T_16959_5 <= _T_9260_3;
              end else begin
                if (_T_10469) begin
                  _T_16959_5 <= _T_9260_4;
                end else begin
                  if (_T_10467) begin
                    _T_16959_5 <= _T_9260_5;
                  end else begin
                    _T_16959_5 <= 8'h0;
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_5 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_6) begin
        if (_T_10499) begin
          _T_16959_6 <= _T_9260_0;
        end else begin
          if (_T_10497) begin
            _T_16959_6 <= _T_9260_1;
          end else begin
            if (_T_10495) begin
              _T_16959_6 <= _T_9260_2;
            end else begin
              if (_T_10493) begin
                _T_16959_6 <= _T_9260_3;
              end else begin
                if (_T_10491) begin
                  _T_16959_6 <= _T_9260_4;
                end else begin
                  if (_T_10489) begin
                    _T_16959_6 <= _T_9260_5;
                  end else begin
                    if (_T_10487) begin
                      _T_16959_6 <= _T_9260_6;
                    end else begin
                      _T_16959_6 <= 8'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_6 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_7) begin
        if (_T_10524) begin
          _T_16959_7 <= _T_9260_0;
        end else begin
          if (_T_10522) begin
            _T_16959_7 <= _T_9260_1;
          end else begin
            if (_T_10520) begin
              _T_16959_7 <= _T_9260_2;
            end else begin
              if (_T_10518) begin
                _T_16959_7 <= _T_9260_3;
              end else begin
                if (_T_10516) begin
                  _T_16959_7 <= _T_9260_4;
                end else begin
                  if (_T_10514) begin
                    _T_16959_7 <= _T_9260_5;
                  end else begin
                    if (_T_10512) begin
                      _T_16959_7 <= _T_9260_6;
                    end else begin
                      if (_T_10510) begin
                        _T_16959_7 <= _T_9260_7;
                      end else begin
                        _T_16959_7 <= 8'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_7 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_8) begin
        if (_T_10552) begin
          _T_16959_8 <= _T_9260_0;
        end else begin
          if (_T_10550) begin
            _T_16959_8 <= _T_9260_1;
          end else begin
            if (_T_10548) begin
              _T_16959_8 <= _T_9260_2;
            end else begin
              if (_T_10546) begin
                _T_16959_8 <= _T_9260_3;
              end else begin
                if (_T_10544) begin
                  _T_16959_8 <= _T_9260_4;
                end else begin
                  if (_T_10542) begin
                    _T_16959_8 <= _T_9260_5;
                  end else begin
                    if (_T_10540) begin
                      _T_16959_8 <= _T_9260_6;
                    end else begin
                      if (_T_10538) begin
                        _T_16959_8 <= _T_9260_7;
                      end else begin
                        if (_T_10536) begin
                          _T_16959_8 <= _T_9260_8;
                        end else begin
                          _T_16959_8 <= 8'h0;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_8 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_9) begin
        if (_T_10583) begin
          _T_16959_9 <= _T_9260_0;
        end else begin
          if (_T_10581) begin
            _T_16959_9 <= _T_9260_1;
          end else begin
            if (_T_10579) begin
              _T_16959_9 <= _T_9260_2;
            end else begin
              if (_T_10577) begin
                _T_16959_9 <= _T_9260_3;
              end else begin
                if (_T_10575) begin
                  _T_16959_9 <= _T_9260_4;
                end else begin
                  if (_T_10573) begin
                    _T_16959_9 <= _T_9260_5;
                  end else begin
                    if (_T_10571) begin
                      _T_16959_9 <= _T_9260_6;
                    end else begin
                      if (_T_10569) begin
                        _T_16959_9 <= _T_9260_7;
                      end else begin
                        if (_T_10567) begin
                          _T_16959_9 <= _T_9260_8;
                        end else begin
                          if (_T_10565) begin
                            _T_16959_9 <= _T_9260_9;
                          end else begin
                            _T_16959_9 <= 8'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_9 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_10) begin
        if (_T_10617) begin
          _T_16959_10 <= _T_9260_0;
        end else begin
          if (_T_10615) begin
            _T_16959_10 <= _T_9260_1;
          end else begin
            if (_T_10613) begin
              _T_16959_10 <= _T_9260_2;
            end else begin
              if (_T_10611) begin
                _T_16959_10 <= _T_9260_3;
              end else begin
                if (_T_10609) begin
                  _T_16959_10 <= _T_9260_4;
                end else begin
                  if (_T_10607) begin
                    _T_16959_10 <= _T_9260_5;
                  end else begin
                    if (_T_10605) begin
                      _T_16959_10 <= _T_9260_6;
                    end else begin
                      if (_T_10603) begin
                        _T_16959_10 <= _T_9260_7;
                      end else begin
                        if (_T_10601) begin
                          _T_16959_10 <= _T_9260_8;
                        end else begin
                          if (_T_10599) begin
                            _T_16959_10 <= _T_9260_9;
                          end else begin
                            if (_T_10597) begin
                              _T_16959_10 <= _T_9260_10;
                            end else begin
                              _T_16959_10 <= 8'h0;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_10 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_11) begin
        if (_T_10654) begin
          _T_16959_11 <= _T_9260_0;
        end else begin
          if (_T_10652) begin
            _T_16959_11 <= _T_9260_1;
          end else begin
            if (_T_10650) begin
              _T_16959_11 <= _T_9260_2;
            end else begin
              if (_T_10648) begin
                _T_16959_11 <= _T_9260_3;
              end else begin
                if (_T_10646) begin
                  _T_16959_11 <= _T_9260_4;
                end else begin
                  if (_T_10644) begin
                    _T_16959_11 <= _T_9260_5;
                  end else begin
                    if (_T_10642) begin
                      _T_16959_11 <= _T_9260_6;
                    end else begin
                      if (_T_10640) begin
                        _T_16959_11 <= _T_9260_7;
                      end else begin
                        if (_T_10638) begin
                          _T_16959_11 <= _T_9260_8;
                        end else begin
                          if (_T_10636) begin
                            _T_16959_11 <= _T_9260_9;
                          end else begin
                            if (_T_10634) begin
                              _T_16959_11 <= _T_9260_10;
                            end else begin
                              if (_T_10632) begin
                                _T_16959_11 <= _T_9260_11;
                              end else begin
                                _T_16959_11 <= 8'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_11 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_12) begin
        if (_T_10694) begin
          _T_16959_12 <= _T_9260_0;
        end else begin
          if (_T_10692) begin
            _T_16959_12 <= _T_9260_1;
          end else begin
            if (_T_10690) begin
              _T_16959_12 <= _T_9260_2;
            end else begin
              if (_T_10688) begin
                _T_16959_12 <= _T_9260_3;
              end else begin
                if (_T_10686) begin
                  _T_16959_12 <= _T_9260_4;
                end else begin
                  if (_T_10684) begin
                    _T_16959_12 <= _T_9260_5;
                  end else begin
                    if (_T_10682) begin
                      _T_16959_12 <= _T_9260_6;
                    end else begin
                      if (_T_10680) begin
                        _T_16959_12 <= _T_9260_7;
                      end else begin
                        if (_T_10678) begin
                          _T_16959_12 <= _T_9260_8;
                        end else begin
                          if (_T_10676) begin
                            _T_16959_12 <= _T_9260_9;
                          end else begin
                            if (_T_10674) begin
                              _T_16959_12 <= _T_9260_10;
                            end else begin
                              if (_T_10672) begin
                                _T_16959_12 <= _T_9260_11;
                              end else begin
                                if (_T_10670) begin
                                  _T_16959_12 <= _T_9260_12;
                                end else begin
                                  _T_16959_12 <= 8'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_12 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_13) begin
        if (_T_10737) begin
          _T_16959_13 <= _T_9260_0;
        end else begin
          if (_T_10735) begin
            _T_16959_13 <= _T_9260_1;
          end else begin
            if (_T_10733) begin
              _T_16959_13 <= _T_9260_2;
            end else begin
              if (_T_10731) begin
                _T_16959_13 <= _T_9260_3;
              end else begin
                if (_T_10729) begin
                  _T_16959_13 <= _T_9260_4;
                end else begin
                  if (_T_10727) begin
                    _T_16959_13 <= _T_9260_5;
                  end else begin
                    if (_T_10725) begin
                      _T_16959_13 <= _T_9260_6;
                    end else begin
                      if (_T_10723) begin
                        _T_16959_13 <= _T_9260_7;
                      end else begin
                        if (_T_10721) begin
                          _T_16959_13 <= _T_9260_8;
                        end else begin
                          if (_T_10719) begin
                            _T_16959_13 <= _T_9260_9;
                          end else begin
                            if (_T_10717) begin
                              _T_16959_13 <= _T_9260_10;
                            end else begin
                              if (_T_10715) begin
                                _T_16959_13 <= _T_9260_11;
                              end else begin
                                if (_T_10713) begin
                                  _T_16959_13 <= _T_9260_12;
                                end else begin
                                  if (_T_10711) begin
                                    _T_16959_13 <= _T_9260_13;
                                  end else begin
                                    _T_16959_13 <= 8'h0;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_13 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_14) begin
        if (_T_10783) begin
          _T_16959_14 <= _T_9260_0;
        end else begin
          if (_T_10781) begin
            _T_16959_14 <= _T_9260_1;
          end else begin
            if (_T_10779) begin
              _T_16959_14 <= _T_9260_2;
            end else begin
              if (_T_10777) begin
                _T_16959_14 <= _T_9260_3;
              end else begin
                if (_T_10775) begin
                  _T_16959_14 <= _T_9260_4;
                end else begin
                  if (_T_10773) begin
                    _T_16959_14 <= _T_9260_5;
                  end else begin
                    if (_T_10771) begin
                      _T_16959_14 <= _T_9260_6;
                    end else begin
                      if (_T_10769) begin
                        _T_16959_14 <= _T_9260_7;
                      end else begin
                        if (_T_10767) begin
                          _T_16959_14 <= _T_9260_8;
                        end else begin
                          if (_T_10765) begin
                            _T_16959_14 <= _T_9260_9;
                          end else begin
                            if (_T_10763) begin
                              _T_16959_14 <= _T_9260_10;
                            end else begin
                              if (_T_10761) begin
                                _T_16959_14 <= _T_9260_11;
                              end else begin
                                if (_T_10759) begin
                                  _T_16959_14 <= _T_9260_12;
                                end else begin
                                  if (_T_10757) begin
                                    _T_16959_14 <= _T_9260_13;
                                  end else begin
                                    if (_T_10755) begin
                                      _T_16959_14 <= _T_9260_14;
                                    end else begin
                                      _T_16959_14 <= 8'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_14 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_15) begin
        if (_T_10832) begin
          _T_16959_15 <= _T_9260_0;
        end else begin
          if (_T_10830) begin
            _T_16959_15 <= _T_9260_1;
          end else begin
            if (_T_10828) begin
              _T_16959_15 <= _T_9260_2;
            end else begin
              if (_T_10826) begin
                _T_16959_15 <= _T_9260_3;
              end else begin
                if (_T_10824) begin
                  _T_16959_15 <= _T_9260_4;
                end else begin
                  if (_T_10822) begin
                    _T_16959_15 <= _T_9260_5;
                  end else begin
                    if (_T_10820) begin
                      _T_16959_15 <= _T_9260_6;
                    end else begin
                      if (_T_10818) begin
                        _T_16959_15 <= _T_9260_7;
                      end else begin
                        if (_T_10816) begin
                          _T_16959_15 <= _T_9260_8;
                        end else begin
                          if (_T_10814) begin
                            _T_16959_15 <= _T_9260_9;
                          end else begin
                            if (_T_10812) begin
                              _T_16959_15 <= _T_9260_10;
                            end else begin
                              if (_T_10810) begin
                                _T_16959_15 <= _T_9260_11;
                              end else begin
                                if (_T_10808) begin
                                  _T_16959_15 <= _T_9260_12;
                                end else begin
                                  if (_T_10806) begin
                                    _T_16959_15 <= _T_9260_13;
                                  end else begin
                                    if (_T_10804) begin
                                      _T_16959_15 <= _T_9260_14;
                                    end else begin
                                      if (_T_10802) begin
                                        _T_16959_15 <= _T_9260_15;
                                      end else begin
                                        _T_16959_15 <= 8'h0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_15 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_16) begin
        if (_T_10884) begin
          _T_16959_16 <= _T_9260_0;
        end else begin
          if (_T_10882) begin
            _T_16959_16 <= _T_9260_1;
          end else begin
            if (_T_10880) begin
              _T_16959_16 <= _T_9260_2;
            end else begin
              if (_T_10878) begin
                _T_16959_16 <= _T_9260_3;
              end else begin
                if (_T_10876) begin
                  _T_16959_16 <= _T_9260_4;
                end else begin
                  if (_T_10874) begin
                    _T_16959_16 <= _T_9260_5;
                  end else begin
                    if (_T_10872) begin
                      _T_16959_16 <= _T_9260_6;
                    end else begin
                      if (_T_10870) begin
                        _T_16959_16 <= _T_9260_7;
                      end else begin
                        if (_T_10868) begin
                          _T_16959_16 <= _T_9260_8;
                        end else begin
                          if (_T_10866) begin
                            _T_16959_16 <= _T_9260_9;
                          end else begin
                            if (_T_10864) begin
                              _T_16959_16 <= _T_9260_10;
                            end else begin
                              if (_T_10862) begin
                                _T_16959_16 <= _T_9260_11;
                              end else begin
                                if (_T_10860) begin
                                  _T_16959_16 <= _T_9260_12;
                                end else begin
                                  if (_T_10858) begin
                                    _T_16959_16 <= _T_9260_13;
                                  end else begin
                                    if (_T_10856) begin
                                      _T_16959_16 <= _T_9260_14;
                                    end else begin
                                      if (_T_10854) begin
                                        _T_16959_16 <= _T_9260_15;
                                      end else begin
                                        if (_T_10852) begin
                                          _T_16959_16 <= _T_9260_16;
                                        end else begin
                                          _T_16959_16 <= 8'h0;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_16 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_17) begin
        if (_T_10939) begin
          _T_16959_17 <= _T_9260_0;
        end else begin
          if (_T_10937) begin
            _T_16959_17 <= _T_9260_1;
          end else begin
            if (_T_10935) begin
              _T_16959_17 <= _T_9260_2;
            end else begin
              if (_T_10933) begin
                _T_16959_17 <= _T_9260_3;
              end else begin
                if (_T_10931) begin
                  _T_16959_17 <= _T_9260_4;
                end else begin
                  if (_T_10929) begin
                    _T_16959_17 <= _T_9260_5;
                  end else begin
                    if (_T_10927) begin
                      _T_16959_17 <= _T_9260_6;
                    end else begin
                      if (_T_10925) begin
                        _T_16959_17 <= _T_9260_7;
                      end else begin
                        if (_T_10923) begin
                          _T_16959_17 <= _T_9260_8;
                        end else begin
                          if (_T_10921) begin
                            _T_16959_17 <= _T_9260_9;
                          end else begin
                            if (_T_10919) begin
                              _T_16959_17 <= _T_9260_10;
                            end else begin
                              if (_T_10917) begin
                                _T_16959_17 <= _T_9260_11;
                              end else begin
                                if (_T_10915) begin
                                  _T_16959_17 <= _T_9260_12;
                                end else begin
                                  if (_T_10913) begin
                                    _T_16959_17 <= _T_9260_13;
                                  end else begin
                                    if (_T_10911) begin
                                      _T_16959_17 <= _T_9260_14;
                                    end else begin
                                      if (_T_10909) begin
                                        _T_16959_17 <= _T_9260_15;
                                      end else begin
                                        if (_T_10907) begin
                                          _T_16959_17 <= _T_9260_16;
                                        end else begin
                                          if (_T_10905) begin
                                            _T_16959_17 <= _T_9260_17;
                                          end else begin
                                            _T_16959_17 <= 8'h0;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_17 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_18) begin
        if (_T_10997) begin
          _T_16959_18 <= _T_9260_0;
        end else begin
          if (_T_10995) begin
            _T_16959_18 <= _T_9260_1;
          end else begin
            if (_T_10993) begin
              _T_16959_18 <= _T_9260_2;
            end else begin
              if (_T_10991) begin
                _T_16959_18 <= _T_9260_3;
              end else begin
                if (_T_10989) begin
                  _T_16959_18 <= _T_9260_4;
                end else begin
                  if (_T_10987) begin
                    _T_16959_18 <= _T_9260_5;
                  end else begin
                    if (_T_10985) begin
                      _T_16959_18 <= _T_9260_6;
                    end else begin
                      if (_T_10983) begin
                        _T_16959_18 <= _T_9260_7;
                      end else begin
                        if (_T_10981) begin
                          _T_16959_18 <= _T_9260_8;
                        end else begin
                          if (_T_10979) begin
                            _T_16959_18 <= _T_9260_9;
                          end else begin
                            if (_T_10977) begin
                              _T_16959_18 <= _T_9260_10;
                            end else begin
                              if (_T_10975) begin
                                _T_16959_18 <= _T_9260_11;
                              end else begin
                                if (_T_10973) begin
                                  _T_16959_18 <= _T_9260_12;
                                end else begin
                                  if (_T_10971) begin
                                    _T_16959_18 <= _T_9260_13;
                                  end else begin
                                    if (_T_10969) begin
                                      _T_16959_18 <= _T_9260_14;
                                    end else begin
                                      if (_T_10967) begin
                                        _T_16959_18 <= _T_9260_15;
                                      end else begin
                                        if (_T_10965) begin
                                          _T_16959_18 <= _T_9260_16;
                                        end else begin
                                          if (_T_10963) begin
                                            _T_16959_18 <= _T_9260_17;
                                          end else begin
                                            if (_T_10961) begin
                                              _T_16959_18 <= _T_9260_18;
                                            end else begin
                                              _T_16959_18 <= 8'h0;
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_18 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_19) begin
        if (_T_11058) begin
          _T_16959_19 <= _T_9260_0;
        end else begin
          if (_T_11056) begin
            _T_16959_19 <= _T_9260_1;
          end else begin
            if (_T_11054) begin
              _T_16959_19 <= _T_9260_2;
            end else begin
              if (_T_11052) begin
                _T_16959_19 <= _T_9260_3;
              end else begin
                if (_T_11050) begin
                  _T_16959_19 <= _T_9260_4;
                end else begin
                  if (_T_11048) begin
                    _T_16959_19 <= _T_9260_5;
                  end else begin
                    if (_T_11046) begin
                      _T_16959_19 <= _T_9260_6;
                    end else begin
                      if (_T_11044) begin
                        _T_16959_19 <= _T_9260_7;
                      end else begin
                        if (_T_11042) begin
                          _T_16959_19 <= _T_9260_8;
                        end else begin
                          if (_T_11040) begin
                            _T_16959_19 <= _T_9260_9;
                          end else begin
                            if (_T_11038) begin
                              _T_16959_19 <= _T_9260_10;
                            end else begin
                              if (_T_11036) begin
                                _T_16959_19 <= _T_9260_11;
                              end else begin
                                if (_T_11034) begin
                                  _T_16959_19 <= _T_9260_12;
                                end else begin
                                  if (_T_11032) begin
                                    _T_16959_19 <= _T_9260_13;
                                  end else begin
                                    if (_T_11030) begin
                                      _T_16959_19 <= _T_9260_14;
                                    end else begin
                                      if (_T_11028) begin
                                        _T_16959_19 <= _T_9260_15;
                                      end else begin
                                        if (_T_11026) begin
                                          _T_16959_19 <= _T_9260_16;
                                        end else begin
                                          if (_T_11024) begin
                                            _T_16959_19 <= _T_9260_17;
                                          end else begin
                                            if (_T_11022) begin
                                              _T_16959_19 <= _T_9260_18;
                                            end else begin
                                              if (_T_11020) begin
                                                _T_16959_19 <= _T_9260_19;
                                              end else begin
                                                _T_16959_19 <= 8'h0;
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_19 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_20) begin
        if (_T_11122) begin
          _T_16959_20 <= _T_9260_0;
        end else begin
          if (_T_11120) begin
            _T_16959_20 <= _T_9260_1;
          end else begin
            if (_T_11118) begin
              _T_16959_20 <= _T_9260_2;
            end else begin
              if (_T_11116) begin
                _T_16959_20 <= _T_9260_3;
              end else begin
                if (_T_11114) begin
                  _T_16959_20 <= _T_9260_4;
                end else begin
                  if (_T_11112) begin
                    _T_16959_20 <= _T_9260_5;
                  end else begin
                    if (_T_11110) begin
                      _T_16959_20 <= _T_9260_6;
                    end else begin
                      if (_T_11108) begin
                        _T_16959_20 <= _T_9260_7;
                      end else begin
                        if (_T_11106) begin
                          _T_16959_20 <= _T_9260_8;
                        end else begin
                          if (_T_11104) begin
                            _T_16959_20 <= _T_9260_9;
                          end else begin
                            if (_T_11102) begin
                              _T_16959_20 <= _T_9260_10;
                            end else begin
                              if (_T_11100) begin
                                _T_16959_20 <= _T_9260_11;
                              end else begin
                                if (_T_11098) begin
                                  _T_16959_20 <= _T_9260_12;
                                end else begin
                                  if (_T_11096) begin
                                    _T_16959_20 <= _T_9260_13;
                                  end else begin
                                    if (_T_11094) begin
                                      _T_16959_20 <= _T_9260_14;
                                    end else begin
                                      if (_T_11092) begin
                                        _T_16959_20 <= _T_9260_15;
                                      end else begin
                                        if (_T_11090) begin
                                          _T_16959_20 <= _T_9260_16;
                                        end else begin
                                          if (_T_11088) begin
                                            _T_16959_20 <= _T_9260_17;
                                          end else begin
                                            if (_T_11086) begin
                                              _T_16959_20 <= _T_9260_18;
                                            end else begin
                                              if (_T_11084) begin
                                                _T_16959_20 <= _T_9260_19;
                                              end else begin
                                                if (_T_11082) begin
                                                  _T_16959_20 <= _T_9260_20;
                                                end else begin
                                                  _T_16959_20 <= 8'h0;
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_20 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_21) begin
        if (_T_11189) begin
          _T_16959_21 <= _T_9260_0;
        end else begin
          if (_T_11187) begin
            _T_16959_21 <= _T_9260_1;
          end else begin
            if (_T_11185) begin
              _T_16959_21 <= _T_9260_2;
            end else begin
              if (_T_11183) begin
                _T_16959_21 <= _T_9260_3;
              end else begin
                if (_T_11181) begin
                  _T_16959_21 <= _T_9260_4;
                end else begin
                  if (_T_11179) begin
                    _T_16959_21 <= _T_9260_5;
                  end else begin
                    if (_T_11177) begin
                      _T_16959_21 <= _T_9260_6;
                    end else begin
                      if (_T_11175) begin
                        _T_16959_21 <= _T_9260_7;
                      end else begin
                        if (_T_11173) begin
                          _T_16959_21 <= _T_9260_8;
                        end else begin
                          if (_T_11171) begin
                            _T_16959_21 <= _T_9260_9;
                          end else begin
                            if (_T_11169) begin
                              _T_16959_21 <= _T_9260_10;
                            end else begin
                              if (_T_11167) begin
                                _T_16959_21 <= _T_9260_11;
                              end else begin
                                if (_T_11165) begin
                                  _T_16959_21 <= _T_9260_12;
                                end else begin
                                  if (_T_11163) begin
                                    _T_16959_21 <= _T_9260_13;
                                  end else begin
                                    if (_T_11161) begin
                                      _T_16959_21 <= _T_9260_14;
                                    end else begin
                                      if (_T_11159) begin
                                        _T_16959_21 <= _T_9260_15;
                                      end else begin
                                        if (_T_11157) begin
                                          _T_16959_21 <= _T_9260_16;
                                        end else begin
                                          if (_T_11155) begin
                                            _T_16959_21 <= _T_9260_17;
                                          end else begin
                                            if (_T_11153) begin
                                              _T_16959_21 <= _T_9260_18;
                                            end else begin
                                              if (_T_11151) begin
                                                _T_16959_21 <= _T_9260_19;
                                              end else begin
                                                if (_T_11149) begin
                                                  _T_16959_21 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11147) begin
                                                    _T_16959_21 <= _T_9260_21;
                                                  end else begin
                                                    _T_16959_21 <= 8'h0;
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_21 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_22) begin
        if (_T_11259) begin
          _T_16959_22 <= _T_9260_0;
        end else begin
          if (_T_11257) begin
            _T_16959_22 <= _T_9260_1;
          end else begin
            if (_T_11255) begin
              _T_16959_22 <= _T_9260_2;
            end else begin
              if (_T_11253) begin
                _T_16959_22 <= _T_9260_3;
              end else begin
                if (_T_11251) begin
                  _T_16959_22 <= _T_9260_4;
                end else begin
                  if (_T_11249) begin
                    _T_16959_22 <= _T_9260_5;
                  end else begin
                    if (_T_11247) begin
                      _T_16959_22 <= _T_9260_6;
                    end else begin
                      if (_T_11245) begin
                        _T_16959_22 <= _T_9260_7;
                      end else begin
                        if (_T_11243) begin
                          _T_16959_22 <= _T_9260_8;
                        end else begin
                          if (_T_11241) begin
                            _T_16959_22 <= _T_9260_9;
                          end else begin
                            if (_T_11239) begin
                              _T_16959_22 <= _T_9260_10;
                            end else begin
                              if (_T_11237) begin
                                _T_16959_22 <= _T_9260_11;
                              end else begin
                                if (_T_11235) begin
                                  _T_16959_22 <= _T_9260_12;
                                end else begin
                                  if (_T_11233) begin
                                    _T_16959_22 <= _T_9260_13;
                                  end else begin
                                    if (_T_11231) begin
                                      _T_16959_22 <= _T_9260_14;
                                    end else begin
                                      if (_T_11229) begin
                                        _T_16959_22 <= _T_9260_15;
                                      end else begin
                                        if (_T_11227) begin
                                          _T_16959_22 <= _T_9260_16;
                                        end else begin
                                          if (_T_11225) begin
                                            _T_16959_22 <= _T_9260_17;
                                          end else begin
                                            if (_T_11223) begin
                                              _T_16959_22 <= _T_9260_18;
                                            end else begin
                                              if (_T_11221) begin
                                                _T_16959_22 <= _T_9260_19;
                                              end else begin
                                                if (_T_11219) begin
                                                  _T_16959_22 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11217) begin
                                                    _T_16959_22 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11215) begin
                                                      _T_16959_22 <= _T_9260_22;
                                                    end else begin
                                                      _T_16959_22 <= 8'h0;
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_22 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_23) begin
        if (_T_11332) begin
          _T_16959_23 <= _T_9260_0;
        end else begin
          if (_T_11330) begin
            _T_16959_23 <= _T_9260_1;
          end else begin
            if (_T_11328) begin
              _T_16959_23 <= _T_9260_2;
            end else begin
              if (_T_11326) begin
                _T_16959_23 <= _T_9260_3;
              end else begin
                if (_T_11324) begin
                  _T_16959_23 <= _T_9260_4;
                end else begin
                  if (_T_11322) begin
                    _T_16959_23 <= _T_9260_5;
                  end else begin
                    if (_T_11320) begin
                      _T_16959_23 <= _T_9260_6;
                    end else begin
                      if (_T_11318) begin
                        _T_16959_23 <= _T_9260_7;
                      end else begin
                        if (_T_11316) begin
                          _T_16959_23 <= _T_9260_8;
                        end else begin
                          if (_T_11314) begin
                            _T_16959_23 <= _T_9260_9;
                          end else begin
                            if (_T_11312) begin
                              _T_16959_23 <= _T_9260_10;
                            end else begin
                              if (_T_11310) begin
                                _T_16959_23 <= _T_9260_11;
                              end else begin
                                if (_T_11308) begin
                                  _T_16959_23 <= _T_9260_12;
                                end else begin
                                  if (_T_11306) begin
                                    _T_16959_23 <= _T_9260_13;
                                  end else begin
                                    if (_T_11304) begin
                                      _T_16959_23 <= _T_9260_14;
                                    end else begin
                                      if (_T_11302) begin
                                        _T_16959_23 <= _T_9260_15;
                                      end else begin
                                        if (_T_11300) begin
                                          _T_16959_23 <= _T_9260_16;
                                        end else begin
                                          if (_T_11298) begin
                                            _T_16959_23 <= _T_9260_17;
                                          end else begin
                                            if (_T_11296) begin
                                              _T_16959_23 <= _T_9260_18;
                                            end else begin
                                              if (_T_11294) begin
                                                _T_16959_23 <= _T_9260_19;
                                              end else begin
                                                if (_T_11292) begin
                                                  _T_16959_23 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11290) begin
                                                    _T_16959_23 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11288) begin
                                                      _T_16959_23 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11286) begin
                                                        _T_16959_23 <= _T_9260_23;
                                                      end else begin
                                                        _T_16959_23 <= 8'h0;
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_23 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_24) begin
        if (_T_11408) begin
          _T_16959_24 <= _T_9260_0;
        end else begin
          if (_T_11406) begin
            _T_16959_24 <= _T_9260_1;
          end else begin
            if (_T_11404) begin
              _T_16959_24 <= _T_9260_2;
            end else begin
              if (_T_11402) begin
                _T_16959_24 <= _T_9260_3;
              end else begin
                if (_T_11400) begin
                  _T_16959_24 <= _T_9260_4;
                end else begin
                  if (_T_11398) begin
                    _T_16959_24 <= _T_9260_5;
                  end else begin
                    if (_T_11396) begin
                      _T_16959_24 <= _T_9260_6;
                    end else begin
                      if (_T_11394) begin
                        _T_16959_24 <= _T_9260_7;
                      end else begin
                        if (_T_11392) begin
                          _T_16959_24 <= _T_9260_8;
                        end else begin
                          if (_T_11390) begin
                            _T_16959_24 <= _T_9260_9;
                          end else begin
                            if (_T_11388) begin
                              _T_16959_24 <= _T_9260_10;
                            end else begin
                              if (_T_11386) begin
                                _T_16959_24 <= _T_9260_11;
                              end else begin
                                if (_T_11384) begin
                                  _T_16959_24 <= _T_9260_12;
                                end else begin
                                  if (_T_11382) begin
                                    _T_16959_24 <= _T_9260_13;
                                  end else begin
                                    if (_T_11380) begin
                                      _T_16959_24 <= _T_9260_14;
                                    end else begin
                                      if (_T_11378) begin
                                        _T_16959_24 <= _T_9260_15;
                                      end else begin
                                        if (_T_11376) begin
                                          _T_16959_24 <= _T_9260_16;
                                        end else begin
                                          if (_T_11374) begin
                                            _T_16959_24 <= _T_9260_17;
                                          end else begin
                                            if (_T_11372) begin
                                              _T_16959_24 <= _T_9260_18;
                                            end else begin
                                              if (_T_11370) begin
                                                _T_16959_24 <= _T_9260_19;
                                              end else begin
                                                if (_T_11368) begin
                                                  _T_16959_24 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11366) begin
                                                    _T_16959_24 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11364) begin
                                                      _T_16959_24 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11362) begin
                                                        _T_16959_24 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11360) begin
                                                          _T_16959_24 <= _T_9260_24;
                                                        end else begin
                                                          _T_16959_24 <= 8'h0;
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_24 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_25) begin
        if (_T_11487) begin
          _T_16959_25 <= _T_9260_0;
        end else begin
          if (_T_11485) begin
            _T_16959_25 <= _T_9260_1;
          end else begin
            if (_T_11483) begin
              _T_16959_25 <= _T_9260_2;
            end else begin
              if (_T_11481) begin
                _T_16959_25 <= _T_9260_3;
              end else begin
                if (_T_11479) begin
                  _T_16959_25 <= _T_9260_4;
                end else begin
                  if (_T_11477) begin
                    _T_16959_25 <= _T_9260_5;
                  end else begin
                    if (_T_11475) begin
                      _T_16959_25 <= _T_9260_6;
                    end else begin
                      if (_T_11473) begin
                        _T_16959_25 <= _T_9260_7;
                      end else begin
                        if (_T_11471) begin
                          _T_16959_25 <= _T_9260_8;
                        end else begin
                          if (_T_11469) begin
                            _T_16959_25 <= _T_9260_9;
                          end else begin
                            if (_T_11467) begin
                              _T_16959_25 <= _T_9260_10;
                            end else begin
                              if (_T_11465) begin
                                _T_16959_25 <= _T_9260_11;
                              end else begin
                                if (_T_11463) begin
                                  _T_16959_25 <= _T_9260_12;
                                end else begin
                                  if (_T_11461) begin
                                    _T_16959_25 <= _T_9260_13;
                                  end else begin
                                    if (_T_11459) begin
                                      _T_16959_25 <= _T_9260_14;
                                    end else begin
                                      if (_T_11457) begin
                                        _T_16959_25 <= _T_9260_15;
                                      end else begin
                                        if (_T_11455) begin
                                          _T_16959_25 <= _T_9260_16;
                                        end else begin
                                          if (_T_11453) begin
                                            _T_16959_25 <= _T_9260_17;
                                          end else begin
                                            if (_T_11451) begin
                                              _T_16959_25 <= _T_9260_18;
                                            end else begin
                                              if (_T_11449) begin
                                                _T_16959_25 <= _T_9260_19;
                                              end else begin
                                                if (_T_11447) begin
                                                  _T_16959_25 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11445) begin
                                                    _T_16959_25 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11443) begin
                                                      _T_16959_25 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11441) begin
                                                        _T_16959_25 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11439) begin
                                                          _T_16959_25 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11437) begin
                                                            _T_16959_25 <= _T_9260_25;
                                                          end else begin
                                                            _T_16959_25 <= 8'h0;
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_25 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_26) begin
        if (_T_11569) begin
          _T_16959_26 <= _T_9260_0;
        end else begin
          if (_T_11567) begin
            _T_16959_26 <= _T_9260_1;
          end else begin
            if (_T_11565) begin
              _T_16959_26 <= _T_9260_2;
            end else begin
              if (_T_11563) begin
                _T_16959_26 <= _T_9260_3;
              end else begin
                if (_T_11561) begin
                  _T_16959_26 <= _T_9260_4;
                end else begin
                  if (_T_11559) begin
                    _T_16959_26 <= _T_9260_5;
                  end else begin
                    if (_T_11557) begin
                      _T_16959_26 <= _T_9260_6;
                    end else begin
                      if (_T_11555) begin
                        _T_16959_26 <= _T_9260_7;
                      end else begin
                        if (_T_11553) begin
                          _T_16959_26 <= _T_9260_8;
                        end else begin
                          if (_T_11551) begin
                            _T_16959_26 <= _T_9260_9;
                          end else begin
                            if (_T_11549) begin
                              _T_16959_26 <= _T_9260_10;
                            end else begin
                              if (_T_11547) begin
                                _T_16959_26 <= _T_9260_11;
                              end else begin
                                if (_T_11545) begin
                                  _T_16959_26 <= _T_9260_12;
                                end else begin
                                  if (_T_11543) begin
                                    _T_16959_26 <= _T_9260_13;
                                  end else begin
                                    if (_T_11541) begin
                                      _T_16959_26 <= _T_9260_14;
                                    end else begin
                                      if (_T_11539) begin
                                        _T_16959_26 <= _T_9260_15;
                                      end else begin
                                        if (_T_11537) begin
                                          _T_16959_26 <= _T_9260_16;
                                        end else begin
                                          if (_T_11535) begin
                                            _T_16959_26 <= _T_9260_17;
                                          end else begin
                                            if (_T_11533) begin
                                              _T_16959_26 <= _T_9260_18;
                                            end else begin
                                              if (_T_11531) begin
                                                _T_16959_26 <= _T_9260_19;
                                              end else begin
                                                if (_T_11529) begin
                                                  _T_16959_26 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11527) begin
                                                    _T_16959_26 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11525) begin
                                                      _T_16959_26 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11523) begin
                                                        _T_16959_26 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11521) begin
                                                          _T_16959_26 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11519) begin
                                                            _T_16959_26 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_11517) begin
                                                              _T_16959_26 <= _T_9260_26;
                                                            end else begin
                                                              _T_16959_26 <= 8'h0;
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_26 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_27) begin
        if (_T_11654) begin
          _T_16959_27 <= _T_9260_0;
        end else begin
          if (_T_11652) begin
            _T_16959_27 <= _T_9260_1;
          end else begin
            if (_T_11650) begin
              _T_16959_27 <= _T_9260_2;
            end else begin
              if (_T_11648) begin
                _T_16959_27 <= _T_9260_3;
              end else begin
                if (_T_11646) begin
                  _T_16959_27 <= _T_9260_4;
                end else begin
                  if (_T_11644) begin
                    _T_16959_27 <= _T_9260_5;
                  end else begin
                    if (_T_11642) begin
                      _T_16959_27 <= _T_9260_6;
                    end else begin
                      if (_T_11640) begin
                        _T_16959_27 <= _T_9260_7;
                      end else begin
                        if (_T_11638) begin
                          _T_16959_27 <= _T_9260_8;
                        end else begin
                          if (_T_11636) begin
                            _T_16959_27 <= _T_9260_9;
                          end else begin
                            if (_T_11634) begin
                              _T_16959_27 <= _T_9260_10;
                            end else begin
                              if (_T_11632) begin
                                _T_16959_27 <= _T_9260_11;
                              end else begin
                                if (_T_11630) begin
                                  _T_16959_27 <= _T_9260_12;
                                end else begin
                                  if (_T_11628) begin
                                    _T_16959_27 <= _T_9260_13;
                                  end else begin
                                    if (_T_11626) begin
                                      _T_16959_27 <= _T_9260_14;
                                    end else begin
                                      if (_T_11624) begin
                                        _T_16959_27 <= _T_9260_15;
                                      end else begin
                                        if (_T_11622) begin
                                          _T_16959_27 <= _T_9260_16;
                                        end else begin
                                          if (_T_11620) begin
                                            _T_16959_27 <= _T_9260_17;
                                          end else begin
                                            if (_T_11618) begin
                                              _T_16959_27 <= _T_9260_18;
                                            end else begin
                                              if (_T_11616) begin
                                                _T_16959_27 <= _T_9260_19;
                                              end else begin
                                                if (_T_11614) begin
                                                  _T_16959_27 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11612) begin
                                                    _T_16959_27 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11610) begin
                                                      _T_16959_27 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11608) begin
                                                        _T_16959_27 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11606) begin
                                                          _T_16959_27 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11604) begin
                                                            _T_16959_27 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_11602) begin
                                                              _T_16959_27 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_11600) begin
                                                                _T_16959_27 <= _T_9260_27;
                                                              end else begin
                                                                _T_16959_27 <= 8'h0;
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_27 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_28) begin
        if (_T_11742) begin
          _T_16959_28 <= _T_9260_0;
        end else begin
          if (_T_11740) begin
            _T_16959_28 <= _T_9260_1;
          end else begin
            if (_T_11738) begin
              _T_16959_28 <= _T_9260_2;
            end else begin
              if (_T_11736) begin
                _T_16959_28 <= _T_9260_3;
              end else begin
                if (_T_11734) begin
                  _T_16959_28 <= _T_9260_4;
                end else begin
                  if (_T_11732) begin
                    _T_16959_28 <= _T_9260_5;
                  end else begin
                    if (_T_11730) begin
                      _T_16959_28 <= _T_9260_6;
                    end else begin
                      if (_T_11728) begin
                        _T_16959_28 <= _T_9260_7;
                      end else begin
                        if (_T_11726) begin
                          _T_16959_28 <= _T_9260_8;
                        end else begin
                          if (_T_11724) begin
                            _T_16959_28 <= _T_9260_9;
                          end else begin
                            if (_T_11722) begin
                              _T_16959_28 <= _T_9260_10;
                            end else begin
                              if (_T_11720) begin
                                _T_16959_28 <= _T_9260_11;
                              end else begin
                                if (_T_11718) begin
                                  _T_16959_28 <= _T_9260_12;
                                end else begin
                                  if (_T_11716) begin
                                    _T_16959_28 <= _T_9260_13;
                                  end else begin
                                    if (_T_11714) begin
                                      _T_16959_28 <= _T_9260_14;
                                    end else begin
                                      if (_T_11712) begin
                                        _T_16959_28 <= _T_9260_15;
                                      end else begin
                                        if (_T_11710) begin
                                          _T_16959_28 <= _T_9260_16;
                                        end else begin
                                          if (_T_11708) begin
                                            _T_16959_28 <= _T_9260_17;
                                          end else begin
                                            if (_T_11706) begin
                                              _T_16959_28 <= _T_9260_18;
                                            end else begin
                                              if (_T_11704) begin
                                                _T_16959_28 <= _T_9260_19;
                                              end else begin
                                                if (_T_11702) begin
                                                  _T_16959_28 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11700) begin
                                                    _T_16959_28 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11698) begin
                                                      _T_16959_28 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11696) begin
                                                        _T_16959_28 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11694) begin
                                                          _T_16959_28 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11692) begin
                                                            _T_16959_28 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_11690) begin
                                                              _T_16959_28 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_11688) begin
                                                                _T_16959_28 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_11686) begin
                                                                  _T_16959_28 <= _T_9260_28;
                                                                end else begin
                                                                  _T_16959_28 <= 8'h0;
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_28 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_29) begin
        if (_T_11833) begin
          _T_16959_29 <= _T_9260_0;
        end else begin
          if (_T_11831) begin
            _T_16959_29 <= _T_9260_1;
          end else begin
            if (_T_11829) begin
              _T_16959_29 <= _T_9260_2;
            end else begin
              if (_T_11827) begin
                _T_16959_29 <= _T_9260_3;
              end else begin
                if (_T_11825) begin
                  _T_16959_29 <= _T_9260_4;
                end else begin
                  if (_T_11823) begin
                    _T_16959_29 <= _T_9260_5;
                  end else begin
                    if (_T_11821) begin
                      _T_16959_29 <= _T_9260_6;
                    end else begin
                      if (_T_11819) begin
                        _T_16959_29 <= _T_9260_7;
                      end else begin
                        if (_T_11817) begin
                          _T_16959_29 <= _T_9260_8;
                        end else begin
                          if (_T_11815) begin
                            _T_16959_29 <= _T_9260_9;
                          end else begin
                            if (_T_11813) begin
                              _T_16959_29 <= _T_9260_10;
                            end else begin
                              if (_T_11811) begin
                                _T_16959_29 <= _T_9260_11;
                              end else begin
                                if (_T_11809) begin
                                  _T_16959_29 <= _T_9260_12;
                                end else begin
                                  if (_T_11807) begin
                                    _T_16959_29 <= _T_9260_13;
                                  end else begin
                                    if (_T_11805) begin
                                      _T_16959_29 <= _T_9260_14;
                                    end else begin
                                      if (_T_11803) begin
                                        _T_16959_29 <= _T_9260_15;
                                      end else begin
                                        if (_T_11801) begin
                                          _T_16959_29 <= _T_9260_16;
                                        end else begin
                                          if (_T_11799) begin
                                            _T_16959_29 <= _T_9260_17;
                                          end else begin
                                            if (_T_11797) begin
                                              _T_16959_29 <= _T_9260_18;
                                            end else begin
                                              if (_T_11795) begin
                                                _T_16959_29 <= _T_9260_19;
                                              end else begin
                                                if (_T_11793) begin
                                                  _T_16959_29 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11791) begin
                                                    _T_16959_29 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11789) begin
                                                      _T_16959_29 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11787) begin
                                                        _T_16959_29 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11785) begin
                                                          _T_16959_29 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11783) begin
                                                            _T_16959_29 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_11781) begin
                                                              _T_16959_29 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_11779) begin
                                                                _T_16959_29 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_11777) begin
                                                                  _T_16959_29 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_11775) begin
                                                                    _T_16959_29 <= _T_9260_29;
                                                                  end else begin
                                                                    _T_16959_29 <= 8'h0;
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_29 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_30) begin
        if (_T_11927) begin
          _T_16959_30 <= _T_9260_0;
        end else begin
          if (_T_11925) begin
            _T_16959_30 <= _T_9260_1;
          end else begin
            if (_T_11923) begin
              _T_16959_30 <= _T_9260_2;
            end else begin
              if (_T_11921) begin
                _T_16959_30 <= _T_9260_3;
              end else begin
                if (_T_11919) begin
                  _T_16959_30 <= _T_9260_4;
                end else begin
                  if (_T_11917) begin
                    _T_16959_30 <= _T_9260_5;
                  end else begin
                    if (_T_11915) begin
                      _T_16959_30 <= _T_9260_6;
                    end else begin
                      if (_T_11913) begin
                        _T_16959_30 <= _T_9260_7;
                      end else begin
                        if (_T_11911) begin
                          _T_16959_30 <= _T_9260_8;
                        end else begin
                          if (_T_11909) begin
                            _T_16959_30 <= _T_9260_9;
                          end else begin
                            if (_T_11907) begin
                              _T_16959_30 <= _T_9260_10;
                            end else begin
                              if (_T_11905) begin
                                _T_16959_30 <= _T_9260_11;
                              end else begin
                                if (_T_11903) begin
                                  _T_16959_30 <= _T_9260_12;
                                end else begin
                                  if (_T_11901) begin
                                    _T_16959_30 <= _T_9260_13;
                                  end else begin
                                    if (_T_11899) begin
                                      _T_16959_30 <= _T_9260_14;
                                    end else begin
                                      if (_T_11897) begin
                                        _T_16959_30 <= _T_9260_15;
                                      end else begin
                                        if (_T_11895) begin
                                          _T_16959_30 <= _T_9260_16;
                                        end else begin
                                          if (_T_11893) begin
                                            _T_16959_30 <= _T_9260_17;
                                          end else begin
                                            if (_T_11891) begin
                                              _T_16959_30 <= _T_9260_18;
                                            end else begin
                                              if (_T_11889) begin
                                                _T_16959_30 <= _T_9260_19;
                                              end else begin
                                                if (_T_11887) begin
                                                  _T_16959_30 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11885) begin
                                                    _T_16959_30 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11883) begin
                                                      _T_16959_30 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11881) begin
                                                        _T_16959_30 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11879) begin
                                                          _T_16959_30 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11877) begin
                                                            _T_16959_30 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_11875) begin
                                                              _T_16959_30 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_11873) begin
                                                                _T_16959_30 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_11871) begin
                                                                  _T_16959_30 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_11869) begin
                                                                    _T_16959_30 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_11867) begin
                                                                      _T_16959_30 <= _T_9260_30;
                                                                    end else begin
                                                                      _T_16959_30 <= 8'h0;
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_30 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_31) begin
        if (_T_12024) begin
          _T_16959_31 <= _T_9260_0;
        end else begin
          if (_T_12022) begin
            _T_16959_31 <= _T_9260_1;
          end else begin
            if (_T_12020) begin
              _T_16959_31 <= _T_9260_2;
            end else begin
              if (_T_12018) begin
                _T_16959_31 <= _T_9260_3;
              end else begin
                if (_T_12016) begin
                  _T_16959_31 <= _T_9260_4;
                end else begin
                  if (_T_12014) begin
                    _T_16959_31 <= _T_9260_5;
                  end else begin
                    if (_T_12012) begin
                      _T_16959_31 <= _T_9260_6;
                    end else begin
                      if (_T_12010) begin
                        _T_16959_31 <= _T_9260_7;
                      end else begin
                        if (_T_12008) begin
                          _T_16959_31 <= _T_9260_8;
                        end else begin
                          if (_T_12006) begin
                            _T_16959_31 <= _T_9260_9;
                          end else begin
                            if (_T_12004) begin
                              _T_16959_31 <= _T_9260_10;
                            end else begin
                              if (_T_12002) begin
                                _T_16959_31 <= _T_9260_11;
                              end else begin
                                if (_T_12000) begin
                                  _T_16959_31 <= _T_9260_12;
                                end else begin
                                  if (_T_11998) begin
                                    _T_16959_31 <= _T_9260_13;
                                  end else begin
                                    if (_T_11996) begin
                                      _T_16959_31 <= _T_9260_14;
                                    end else begin
                                      if (_T_11994) begin
                                        _T_16959_31 <= _T_9260_15;
                                      end else begin
                                        if (_T_11992) begin
                                          _T_16959_31 <= _T_9260_16;
                                        end else begin
                                          if (_T_11990) begin
                                            _T_16959_31 <= _T_9260_17;
                                          end else begin
                                            if (_T_11988) begin
                                              _T_16959_31 <= _T_9260_18;
                                            end else begin
                                              if (_T_11986) begin
                                                _T_16959_31 <= _T_9260_19;
                                              end else begin
                                                if (_T_11984) begin
                                                  _T_16959_31 <= _T_9260_20;
                                                end else begin
                                                  if (_T_11982) begin
                                                    _T_16959_31 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_11980) begin
                                                      _T_16959_31 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_11978) begin
                                                        _T_16959_31 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_11976) begin
                                                          _T_16959_31 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_11974) begin
                                                            _T_16959_31 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_11972) begin
                                                              _T_16959_31 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_11970) begin
                                                                _T_16959_31 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_11968) begin
                                                                  _T_16959_31 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_11966) begin
                                                                    _T_16959_31 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_11964) begin
                                                                      _T_16959_31 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_11962) begin
                                                                        _T_16959_31 <= _T_9260_31;
                                                                      end else begin
                                                                        _T_16959_31 <= 8'h0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_31 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_32) begin
        if (_T_12124) begin
          _T_16959_32 <= _T_9260_0;
        end else begin
          if (_T_12122) begin
            _T_16959_32 <= _T_9260_1;
          end else begin
            if (_T_12120) begin
              _T_16959_32 <= _T_9260_2;
            end else begin
              if (_T_12118) begin
                _T_16959_32 <= _T_9260_3;
              end else begin
                if (_T_12116) begin
                  _T_16959_32 <= _T_9260_4;
                end else begin
                  if (_T_12114) begin
                    _T_16959_32 <= _T_9260_5;
                  end else begin
                    if (_T_12112) begin
                      _T_16959_32 <= _T_9260_6;
                    end else begin
                      if (_T_12110) begin
                        _T_16959_32 <= _T_9260_7;
                      end else begin
                        if (_T_12108) begin
                          _T_16959_32 <= _T_9260_8;
                        end else begin
                          if (_T_12106) begin
                            _T_16959_32 <= _T_9260_9;
                          end else begin
                            if (_T_12104) begin
                              _T_16959_32 <= _T_9260_10;
                            end else begin
                              if (_T_12102) begin
                                _T_16959_32 <= _T_9260_11;
                              end else begin
                                if (_T_12100) begin
                                  _T_16959_32 <= _T_9260_12;
                                end else begin
                                  if (_T_12098) begin
                                    _T_16959_32 <= _T_9260_13;
                                  end else begin
                                    if (_T_12096) begin
                                      _T_16959_32 <= _T_9260_14;
                                    end else begin
                                      if (_T_12094) begin
                                        _T_16959_32 <= _T_9260_15;
                                      end else begin
                                        if (_T_12092) begin
                                          _T_16959_32 <= _T_9260_16;
                                        end else begin
                                          if (_T_12090) begin
                                            _T_16959_32 <= _T_9260_17;
                                          end else begin
                                            if (_T_12088) begin
                                              _T_16959_32 <= _T_9260_18;
                                            end else begin
                                              if (_T_12086) begin
                                                _T_16959_32 <= _T_9260_19;
                                              end else begin
                                                if (_T_12084) begin
                                                  _T_16959_32 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12082) begin
                                                    _T_16959_32 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12080) begin
                                                      _T_16959_32 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12078) begin
                                                        _T_16959_32 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12076) begin
                                                          _T_16959_32 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12074) begin
                                                            _T_16959_32 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12072) begin
                                                              _T_16959_32 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12070) begin
                                                                _T_16959_32 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12068) begin
                                                                  _T_16959_32 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12066) begin
                                                                    _T_16959_32 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12064) begin
                                                                      _T_16959_32 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12062) begin
                                                                        _T_16959_32 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12060) begin
                                                                          _T_16959_32 <= _T_9260_32;
                                                                        end else begin
                                                                          _T_16959_32 <= 8'h0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_32 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_33) begin
        if (_T_12227) begin
          _T_16959_33 <= _T_9260_0;
        end else begin
          if (_T_12225) begin
            _T_16959_33 <= _T_9260_1;
          end else begin
            if (_T_12223) begin
              _T_16959_33 <= _T_9260_2;
            end else begin
              if (_T_12221) begin
                _T_16959_33 <= _T_9260_3;
              end else begin
                if (_T_12219) begin
                  _T_16959_33 <= _T_9260_4;
                end else begin
                  if (_T_12217) begin
                    _T_16959_33 <= _T_9260_5;
                  end else begin
                    if (_T_12215) begin
                      _T_16959_33 <= _T_9260_6;
                    end else begin
                      if (_T_12213) begin
                        _T_16959_33 <= _T_9260_7;
                      end else begin
                        if (_T_12211) begin
                          _T_16959_33 <= _T_9260_8;
                        end else begin
                          if (_T_12209) begin
                            _T_16959_33 <= _T_9260_9;
                          end else begin
                            if (_T_12207) begin
                              _T_16959_33 <= _T_9260_10;
                            end else begin
                              if (_T_12205) begin
                                _T_16959_33 <= _T_9260_11;
                              end else begin
                                if (_T_12203) begin
                                  _T_16959_33 <= _T_9260_12;
                                end else begin
                                  if (_T_12201) begin
                                    _T_16959_33 <= _T_9260_13;
                                  end else begin
                                    if (_T_12199) begin
                                      _T_16959_33 <= _T_9260_14;
                                    end else begin
                                      if (_T_12197) begin
                                        _T_16959_33 <= _T_9260_15;
                                      end else begin
                                        if (_T_12195) begin
                                          _T_16959_33 <= _T_9260_16;
                                        end else begin
                                          if (_T_12193) begin
                                            _T_16959_33 <= _T_9260_17;
                                          end else begin
                                            if (_T_12191) begin
                                              _T_16959_33 <= _T_9260_18;
                                            end else begin
                                              if (_T_12189) begin
                                                _T_16959_33 <= _T_9260_19;
                                              end else begin
                                                if (_T_12187) begin
                                                  _T_16959_33 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12185) begin
                                                    _T_16959_33 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12183) begin
                                                      _T_16959_33 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12181) begin
                                                        _T_16959_33 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12179) begin
                                                          _T_16959_33 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12177) begin
                                                            _T_16959_33 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12175) begin
                                                              _T_16959_33 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12173) begin
                                                                _T_16959_33 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12171) begin
                                                                  _T_16959_33 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12169) begin
                                                                    _T_16959_33 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12167) begin
                                                                      _T_16959_33 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12165) begin
                                                                        _T_16959_33 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12163) begin
                                                                          _T_16959_33 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12161) begin
                                                                            _T_16959_33 <= _T_9260_33;
                                                                          end else begin
                                                                            _T_16959_33 <= 8'h0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_33 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_34) begin
        if (_T_12333) begin
          _T_16959_34 <= _T_9260_0;
        end else begin
          if (_T_12331) begin
            _T_16959_34 <= _T_9260_1;
          end else begin
            if (_T_12329) begin
              _T_16959_34 <= _T_9260_2;
            end else begin
              if (_T_12327) begin
                _T_16959_34 <= _T_9260_3;
              end else begin
                if (_T_12325) begin
                  _T_16959_34 <= _T_9260_4;
                end else begin
                  if (_T_12323) begin
                    _T_16959_34 <= _T_9260_5;
                  end else begin
                    if (_T_12321) begin
                      _T_16959_34 <= _T_9260_6;
                    end else begin
                      if (_T_12319) begin
                        _T_16959_34 <= _T_9260_7;
                      end else begin
                        if (_T_12317) begin
                          _T_16959_34 <= _T_9260_8;
                        end else begin
                          if (_T_12315) begin
                            _T_16959_34 <= _T_9260_9;
                          end else begin
                            if (_T_12313) begin
                              _T_16959_34 <= _T_9260_10;
                            end else begin
                              if (_T_12311) begin
                                _T_16959_34 <= _T_9260_11;
                              end else begin
                                if (_T_12309) begin
                                  _T_16959_34 <= _T_9260_12;
                                end else begin
                                  if (_T_12307) begin
                                    _T_16959_34 <= _T_9260_13;
                                  end else begin
                                    if (_T_12305) begin
                                      _T_16959_34 <= _T_9260_14;
                                    end else begin
                                      if (_T_12303) begin
                                        _T_16959_34 <= _T_9260_15;
                                      end else begin
                                        if (_T_12301) begin
                                          _T_16959_34 <= _T_9260_16;
                                        end else begin
                                          if (_T_12299) begin
                                            _T_16959_34 <= _T_9260_17;
                                          end else begin
                                            if (_T_12297) begin
                                              _T_16959_34 <= _T_9260_18;
                                            end else begin
                                              if (_T_12295) begin
                                                _T_16959_34 <= _T_9260_19;
                                              end else begin
                                                if (_T_12293) begin
                                                  _T_16959_34 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12291) begin
                                                    _T_16959_34 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12289) begin
                                                      _T_16959_34 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12287) begin
                                                        _T_16959_34 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12285) begin
                                                          _T_16959_34 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12283) begin
                                                            _T_16959_34 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12281) begin
                                                              _T_16959_34 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12279) begin
                                                                _T_16959_34 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12277) begin
                                                                  _T_16959_34 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12275) begin
                                                                    _T_16959_34 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12273) begin
                                                                      _T_16959_34 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12271) begin
                                                                        _T_16959_34 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12269) begin
                                                                          _T_16959_34 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12267) begin
                                                                            _T_16959_34 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12265) begin
                                                                              _T_16959_34 <= _T_9260_34;
                                                                            end else begin
                                                                              _T_16959_34 <= 8'h0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_34 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_35) begin
        if (_T_12442) begin
          _T_16959_35 <= _T_9260_0;
        end else begin
          if (_T_12440) begin
            _T_16959_35 <= _T_9260_1;
          end else begin
            if (_T_12438) begin
              _T_16959_35 <= _T_9260_2;
            end else begin
              if (_T_12436) begin
                _T_16959_35 <= _T_9260_3;
              end else begin
                if (_T_12434) begin
                  _T_16959_35 <= _T_9260_4;
                end else begin
                  if (_T_12432) begin
                    _T_16959_35 <= _T_9260_5;
                  end else begin
                    if (_T_12430) begin
                      _T_16959_35 <= _T_9260_6;
                    end else begin
                      if (_T_12428) begin
                        _T_16959_35 <= _T_9260_7;
                      end else begin
                        if (_T_12426) begin
                          _T_16959_35 <= _T_9260_8;
                        end else begin
                          if (_T_12424) begin
                            _T_16959_35 <= _T_9260_9;
                          end else begin
                            if (_T_12422) begin
                              _T_16959_35 <= _T_9260_10;
                            end else begin
                              if (_T_12420) begin
                                _T_16959_35 <= _T_9260_11;
                              end else begin
                                if (_T_12418) begin
                                  _T_16959_35 <= _T_9260_12;
                                end else begin
                                  if (_T_12416) begin
                                    _T_16959_35 <= _T_9260_13;
                                  end else begin
                                    if (_T_12414) begin
                                      _T_16959_35 <= _T_9260_14;
                                    end else begin
                                      if (_T_12412) begin
                                        _T_16959_35 <= _T_9260_15;
                                      end else begin
                                        if (_T_12410) begin
                                          _T_16959_35 <= _T_9260_16;
                                        end else begin
                                          if (_T_12408) begin
                                            _T_16959_35 <= _T_9260_17;
                                          end else begin
                                            if (_T_12406) begin
                                              _T_16959_35 <= _T_9260_18;
                                            end else begin
                                              if (_T_12404) begin
                                                _T_16959_35 <= _T_9260_19;
                                              end else begin
                                                if (_T_12402) begin
                                                  _T_16959_35 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12400) begin
                                                    _T_16959_35 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12398) begin
                                                      _T_16959_35 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12396) begin
                                                        _T_16959_35 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12394) begin
                                                          _T_16959_35 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12392) begin
                                                            _T_16959_35 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12390) begin
                                                              _T_16959_35 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12388) begin
                                                                _T_16959_35 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12386) begin
                                                                  _T_16959_35 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12384) begin
                                                                    _T_16959_35 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12382) begin
                                                                      _T_16959_35 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12380) begin
                                                                        _T_16959_35 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12378) begin
                                                                          _T_16959_35 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12376) begin
                                                                            _T_16959_35 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12374) begin
                                                                              _T_16959_35 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_12372) begin
                                                                                _T_16959_35 <= _T_9260_35;
                                                                              end else begin
                                                                                _T_16959_35 <= 8'h0;
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_35 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_36) begin
        if (_T_12554) begin
          _T_16959_36 <= _T_9260_0;
        end else begin
          if (_T_12552) begin
            _T_16959_36 <= _T_9260_1;
          end else begin
            if (_T_12550) begin
              _T_16959_36 <= _T_9260_2;
            end else begin
              if (_T_12548) begin
                _T_16959_36 <= _T_9260_3;
              end else begin
                if (_T_12546) begin
                  _T_16959_36 <= _T_9260_4;
                end else begin
                  if (_T_12544) begin
                    _T_16959_36 <= _T_9260_5;
                  end else begin
                    if (_T_12542) begin
                      _T_16959_36 <= _T_9260_6;
                    end else begin
                      if (_T_12540) begin
                        _T_16959_36 <= _T_9260_7;
                      end else begin
                        if (_T_12538) begin
                          _T_16959_36 <= _T_9260_8;
                        end else begin
                          if (_T_12536) begin
                            _T_16959_36 <= _T_9260_9;
                          end else begin
                            if (_T_12534) begin
                              _T_16959_36 <= _T_9260_10;
                            end else begin
                              if (_T_12532) begin
                                _T_16959_36 <= _T_9260_11;
                              end else begin
                                if (_T_12530) begin
                                  _T_16959_36 <= _T_9260_12;
                                end else begin
                                  if (_T_12528) begin
                                    _T_16959_36 <= _T_9260_13;
                                  end else begin
                                    if (_T_12526) begin
                                      _T_16959_36 <= _T_9260_14;
                                    end else begin
                                      if (_T_12524) begin
                                        _T_16959_36 <= _T_9260_15;
                                      end else begin
                                        if (_T_12522) begin
                                          _T_16959_36 <= _T_9260_16;
                                        end else begin
                                          if (_T_12520) begin
                                            _T_16959_36 <= _T_9260_17;
                                          end else begin
                                            if (_T_12518) begin
                                              _T_16959_36 <= _T_9260_18;
                                            end else begin
                                              if (_T_12516) begin
                                                _T_16959_36 <= _T_9260_19;
                                              end else begin
                                                if (_T_12514) begin
                                                  _T_16959_36 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12512) begin
                                                    _T_16959_36 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12510) begin
                                                      _T_16959_36 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12508) begin
                                                        _T_16959_36 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12506) begin
                                                          _T_16959_36 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12504) begin
                                                            _T_16959_36 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12502) begin
                                                              _T_16959_36 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12500) begin
                                                                _T_16959_36 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12498) begin
                                                                  _T_16959_36 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12496) begin
                                                                    _T_16959_36 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12494) begin
                                                                      _T_16959_36 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12492) begin
                                                                        _T_16959_36 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12490) begin
                                                                          _T_16959_36 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12488) begin
                                                                            _T_16959_36 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12486) begin
                                                                              _T_16959_36 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_12484) begin
                                                                                _T_16959_36 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_12482) begin
                                                                                  _T_16959_36 <= _T_9260_36;
                                                                                end else begin
                                                                                  _T_16959_36 <= 8'h0;
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_36 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_37) begin
        if (_T_12669) begin
          _T_16959_37 <= _T_9260_0;
        end else begin
          if (_T_12667) begin
            _T_16959_37 <= _T_9260_1;
          end else begin
            if (_T_12665) begin
              _T_16959_37 <= _T_9260_2;
            end else begin
              if (_T_12663) begin
                _T_16959_37 <= _T_9260_3;
              end else begin
                if (_T_12661) begin
                  _T_16959_37 <= _T_9260_4;
                end else begin
                  if (_T_12659) begin
                    _T_16959_37 <= _T_9260_5;
                  end else begin
                    if (_T_12657) begin
                      _T_16959_37 <= _T_9260_6;
                    end else begin
                      if (_T_12655) begin
                        _T_16959_37 <= _T_9260_7;
                      end else begin
                        if (_T_12653) begin
                          _T_16959_37 <= _T_9260_8;
                        end else begin
                          if (_T_12651) begin
                            _T_16959_37 <= _T_9260_9;
                          end else begin
                            if (_T_12649) begin
                              _T_16959_37 <= _T_9260_10;
                            end else begin
                              if (_T_12647) begin
                                _T_16959_37 <= _T_9260_11;
                              end else begin
                                if (_T_12645) begin
                                  _T_16959_37 <= _T_9260_12;
                                end else begin
                                  if (_T_12643) begin
                                    _T_16959_37 <= _T_9260_13;
                                  end else begin
                                    if (_T_12641) begin
                                      _T_16959_37 <= _T_9260_14;
                                    end else begin
                                      if (_T_12639) begin
                                        _T_16959_37 <= _T_9260_15;
                                      end else begin
                                        if (_T_12637) begin
                                          _T_16959_37 <= _T_9260_16;
                                        end else begin
                                          if (_T_12635) begin
                                            _T_16959_37 <= _T_9260_17;
                                          end else begin
                                            if (_T_12633) begin
                                              _T_16959_37 <= _T_9260_18;
                                            end else begin
                                              if (_T_12631) begin
                                                _T_16959_37 <= _T_9260_19;
                                              end else begin
                                                if (_T_12629) begin
                                                  _T_16959_37 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12627) begin
                                                    _T_16959_37 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12625) begin
                                                      _T_16959_37 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12623) begin
                                                        _T_16959_37 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12621) begin
                                                          _T_16959_37 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12619) begin
                                                            _T_16959_37 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12617) begin
                                                              _T_16959_37 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12615) begin
                                                                _T_16959_37 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12613) begin
                                                                  _T_16959_37 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12611) begin
                                                                    _T_16959_37 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12609) begin
                                                                      _T_16959_37 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12607) begin
                                                                        _T_16959_37 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12605) begin
                                                                          _T_16959_37 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12603) begin
                                                                            _T_16959_37 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12601) begin
                                                                              _T_16959_37 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_12599) begin
                                                                                _T_16959_37 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_12597) begin
                                                                                  _T_16959_37 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_12595) begin
                                                                                    _T_16959_37 <= _T_9260_37;
                                                                                  end else begin
                                                                                    _T_16959_37 <= 8'h0;
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_37 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_38) begin
        if (_T_12787) begin
          _T_16959_38 <= _T_9260_0;
        end else begin
          if (_T_12785) begin
            _T_16959_38 <= _T_9260_1;
          end else begin
            if (_T_12783) begin
              _T_16959_38 <= _T_9260_2;
            end else begin
              if (_T_12781) begin
                _T_16959_38 <= _T_9260_3;
              end else begin
                if (_T_12779) begin
                  _T_16959_38 <= _T_9260_4;
                end else begin
                  if (_T_12777) begin
                    _T_16959_38 <= _T_9260_5;
                  end else begin
                    if (_T_12775) begin
                      _T_16959_38 <= _T_9260_6;
                    end else begin
                      if (_T_12773) begin
                        _T_16959_38 <= _T_9260_7;
                      end else begin
                        if (_T_12771) begin
                          _T_16959_38 <= _T_9260_8;
                        end else begin
                          if (_T_12769) begin
                            _T_16959_38 <= _T_9260_9;
                          end else begin
                            if (_T_12767) begin
                              _T_16959_38 <= _T_9260_10;
                            end else begin
                              if (_T_12765) begin
                                _T_16959_38 <= _T_9260_11;
                              end else begin
                                if (_T_12763) begin
                                  _T_16959_38 <= _T_9260_12;
                                end else begin
                                  if (_T_12761) begin
                                    _T_16959_38 <= _T_9260_13;
                                  end else begin
                                    if (_T_12759) begin
                                      _T_16959_38 <= _T_9260_14;
                                    end else begin
                                      if (_T_12757) begin
                                        _T_16959_38 <= _T_9260_15;
                                      end else begin
                                        if (_T_12755) begin
                                          _T_16959_38 <= _T_9260_16;
                                        end else begin
                                          if (_T_12753) begin
                                            _T_16959_38 <= _T_9260_17;
                                          end else begin
                                            if (_T_12751) begin
                                              _T_16959_38 <= _T_9260_18;
                                            end else begin
                                              if (_T_12749) begin
                                                _T_16959_38 <= _T_9260_19;
                                              end else begin
                                                if (_T_12747) begin
                                                  _T_16959_38 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12745) begin
                                                    _T_16959_38 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12743) begin
                                                      _T_16959_38 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12741) begin
                                                        _T_16959_38 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12739) begin
                                                          _T_16959_38 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12737) begin
                                                            _T_16959_38 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12735) begin
                                                              _T_16959_38 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12733) begin
                                                                _T_16959_38 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12731) begin
                                                                  _T_16959_38 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12729) begin
                                                                    _T_16959_38 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12727) begin
                                                                      _T_16959_38 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12725) begin
                                                                        _T_16959_38 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12723) begin
                                                                          _T_16959_38 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12721) begin
                                                                            _T_16959_38 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12719) begin
                                                                              _T_16959_38 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_12717) begin
                                                                                _T_16959_38 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_12715) begin
                                                                                  _T_16959_38 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_12713) begin
                                                                                    _T_16959_38 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_12711) begin
                                                                                      _T_16959_38 <= _T_9260_38;
                                                                                    end else begin
                                                                                      _T_16959_38 <= 8'h0;
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_38 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_39) begin
        if (_T_12908) begin
          _T_16959_39 <= _T_9260_0;
        end else begin
          if (_T_12906) begin
            _T_16959_39 <= _T_9260_1;
          end else begin
            if (_T_12904) begin
              _T_16959_39 <= _T_9260_2;
            end else begin
              if (_T_12902) begin
                _T_16959_39 <= _T_9260_3;
              end else begin
                if (_T_12900) begin
                  _T_16959_39 <= _T_9260_4;
                end else begin
                  if (_T_12898) begin
                    _T_16959_39 <= _T_9260_5;
                  end else begin
                    if (_T_12896) begin
                      _T_16959_39 <= _T_9260_6;
                    end else begin
                      if (_T_12894) begin
                        _T_16959_39 <= _T_9260_7;
                      end else begin
                        if (_T_12892) begin
                          _T_16959_39 <= _T_9260_8;
                        end else begin
                          if (_T_12890) begin
                            _T_16959_39 <= _T_9260_9;
                          end else begin
                            if (_T_12888) begin
                              _T_16959_39 <= _T_9260_10;
                            end else begin
                              if (_T_12886) begin
                                _T_16959_39 <= _T_9260_11;
                              end else begin
                                if (_T_12884) begin
                                  _T_16959_39 <= _T_9260_12;
                                end else begin
                                  if (_T_12882) begin
                                    _T_16959_39 <= _T_9260_13;
                                  end else begin
                                    if (_T_12880) begin
                                      _T_16959_39 <= _T_9260_14;
                                    end else begin
                                      if (_T_12878) begin
                                        _T_16959_39 <= _T_9260_15;
                                      end else begin
                                        if (_T_12876) begin
                                          _T_16959_39 <= _T_9260_16;
                                        end else begin
                                          if (_T_12874) begin
                                            _T_16959_39 <= _T_9260_17;
                                          end else begin
                                            if (_T_12872) begin
                                              _T_16959_39 <= _T_9260_18;
                                            end else begin
                                              if (_T_12870) begin
                                                _T_16959_39 <= _T_9260_19;
                                              end else begin
                                                if (_T_12868) begin
                                                  _T_16959_39 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12866) begin
                                                    _T_16959_39 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12864) begin
                                                      _T_16959_39 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12862) begin
                                                        _T_16959_39 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12860) begin
                                                          _T_16959_39 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12858) begin
                                                            _T_16959_39 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12856) begin
                                                              _T_16959_39 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12854) begin
                                                                _T_16959_39 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12852) begin
                                                                  _T_16959_39 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12850) begin
                                                                    _T_16959_39 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12848) begin
                                                                      _T_16959_39 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12846) begin
                                                                        _T_16959_39 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12844) begin
                                                                          _T_16959_39 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12842) begin
                                                                            _T_16959_39 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12840) begin
                                                                              _T_16959_39 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_12838) begin
                                                                                _T_16959_39 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_12836) begin
                                                                                  _T_16959_39 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_12834) begin
                                                                                    _T_16959_39 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_12832) begin
                                                                                      _T_16959_39 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_12830) begin
                                                                                        _T_16959_39 <= _T_9260_39;
                                                                                      end else begin
                                                                                        _T_16959_39 <= 8'h0;
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_39 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_40) begin
        if (_T_13032) begin
          _T_16959_40 <= _T_9260_0;
        end else begin
          if (_T_13030) begin
            _T_16959_40 <= _T_9260_1;
          end else begin
            if (_T_13028) begin
              _T_16959_40 <= _T_9260_2;
            end else begin
              if (_T_13026) begin
                _T_16959_40 <= _T_9260_3;
              end else begin
                if (_T_13024) begin
                  _T_16959_40 <= _T_9260_4;
                end else begin
                  if (_T_13022) begin
                    _T_16959_40 <= _T_9260_5;
                  end else begin
                    if (_T_13020) begin
                      _T_16959_40 <= _T_9260_6;
                    end else begin
                      if (_T_13018) begin
                        _T_16959_40 <= _T_9260_7;
                      end else begin
                        if (_T_13016) begin
                          _T_16959_40 <= _T_9260_8;
                        end else begin
                          if (_T_13014) begin
                            _T_16959_40 <= _T_9260_9;
                          end else begin
                            if (_T_13012) begin
                              _T_16959_40 <= _T_9260_10;
                            end else begin
                              if (_T_13010) begin
                                _T_16959_40 <= _T_9260_11;
                              end else begin
                                if (_T_13008) begin
                                  _T_16959_40 <= _T_9260_12;
                                end else begin
                                  if (_T_13006) begin
                                    _T_16959_40 <= _T_9260_13;
                                  end else begin
                                    if (_T_13004) begin
                                      _T_16959_40 <= _T_9260_14;
                                    end else begin
                                      if (_T_13002) begin
                                        _T_16959_40 <= _T_9260_15;
                                      end else begin
                                        if (_T_13000) begin
                                          _T_16959_40 <= _T_9260_16;
                                        end else begin
                                          if (_T_12998) begin
                                            _T_16959_40 <= _T_9260_17;
                                          end else begin
                                            if (_T_12996) begin
                                              _T_16959_40 <= _T_9260_18;
                                            end else begin
                                              if (_T_12994) begin
                                                _T_16959_40 <= _T_9260_19;
                                              end else begin
                                                if (_T_12992) begin
                                                  _T_16959_40 <= _T_9260_20;
                                                end else begin
                                                  if (_T_12990) begin
                                                    _T_16959_40 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_12988) begin
                                                      _T_16959_40 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_12986) begin
                                                        _T_16959_40 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_12984) begin
                                                          _T_16959_40 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_12982) begin
                                                            _T_16959_40 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_12980) begin
                                                              _T_16959_40 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_12978) begin
                                                                _T_16959_40 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_12976) begin
                                                                  _T_16959_40 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_12974) begin
                                                                    _T_16959_40 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_12972) begin
                                                                      _T_16959_40 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_12970) begin
                                                                        _T_16959_40 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_12968) begin
                                                                          _T_16959_40 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_12966) begin
                                                                            _T_16959_40 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_12964) begin
                                                                              _T_16959_40 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_12962) begin
                                                                                _T_16959_40 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_12960) begin
                                                                                  _T_16959_40 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_12958) begin
                                                                                    _T_16959_40 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_12956) begin
                                                                                      _T_16959_40 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_12954) begin
                                                                                        _T_16959_40 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_12952) begin
                                                                                          _T_16959_40 <= _T_9260_40;
                                                                                        end else begin
                                                                                          _T_16959_40 <= 8'h0;
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_40 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_41) begin
        if (_T_13159) begin
          _T_16959_41 <= _T_9260_0;
        end else begin
          if (_T_13157) begin
            _T_16959_41 <= _T_9260_1;
          end else begin
            if (_T_13155) begin
              _T_16959_41 <= _T_9260_2;
            end else begin
              if (_T_13153) begin
                _T_16959_41 <= _T_9260_3;
              end else begin
                if (_T_13151) begin
                  _T_16959_41 <= _T_9260_4;
                end else begin
                  if (_T_13149) begin
                    _T_16959_41 <= _T_9260_5;
                  end else begin
                    if (_T_13147) begin
                      _T_16959_41 <= _T_9260_6;
                    end else begin
                      if (_T_13145) begin
                        _T_16959_41 <= _T_9260_7;
                      end else begin
                        if (_T_13143) begin
                          _T_16959_41 <= _T_9260_8;
                        end else begin
                          if (_T_13141) begin
                            _T_16959_41 <= _T_9260_9;
                          end else begin
                            if (_T_13139) begin
                              _T_16959_41 <= _T_9260_10;
                            end else begin
                              if (_T_13137) begin
                                _T_16959_41 <= _T_9260_11;
                              end else begin
                                if (_T_13135) begin
                                  _T_16959_41 <= _T_9260_12;
                                end else begin
                                  if (_T_13133) begin
                                    _T_16959_41 <= _T_9260_13;
                                  end else begin
                                    if (_T_13131) begin
                                      _T_16959_41 <= _T_9260_14;
                                    end else begin
                                      if (_T_13129) begin
                                        _T_16959_41 <= _T_9260_15;
                                      end else begin
                                        if (_T_13127) begin
                                          _T_16959_41 <= _T_9260_16;
                                        end else begin
                                          if (_T_13125) begin
                                            _T_16959_41 <= _T_9260_17;
                                          end else begin
                                            if (_T_13123) begin
                                              _T_16959_41 <= _T_9260_18;
                                            end else begin
                                              if (_T_13121) begin
                                                _T_16959_41 <= _T_9260_19;
                                              end else begin
                                                if (_T_13119) begin
                                                  _T_16959_41 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13117) begin
                                                    _T_16959_41 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13115) begin
                                                      _T_16959_41 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13113) begin
                                                        _T_16959_41 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13111) begin
                                                          _T_16959_41 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13109) begin
                                                            _T_16959_41 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13107) begin
                                                              _T_16959_41 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13105) begin
                                                                _T_16959_41 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13103) begin
                                                                  _T_16959_41 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13101) begin
                                                                    _T_16959_41 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13099) begin
                                                                      _T_16959_41 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13097) begin
                                                                        _T_16959_41 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13095) begin
                                                                          _T_16959_41 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13093) begin
                                                                            _T_16959_41 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13091) begin
                                                                              _T_16959_41 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13089) begin
                                                                                _T_16959_41 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13087) begin
                                                                                  _T_16959_41 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13085) begin
                                                                                    _T_16959_41 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13083) begin
                                                                                      _T_16959_41 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13081) begin
                                                                                        _T_16959_41 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13079) begin
                                                                                          _T_16959_41 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13077) begin
                                                                                            _T_16959_41 <= _T_9260_41;
                                                                                          end else begin
                                                                                            _T_16959_41 <= 8'h0;
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_41 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_42) begin
        if (_T_13289) begin
          _T_16959_42 <= _T_9260_0;
        end else begin
          if (_T_13287) begin
            _T_16959_42 <= _T_9260_1;
          end else begin
            if (_T_13285) begin
              _T_16959_42 <= _T_9260_2;
            end else begin
              if (_T_13283) begin
                _T_16959_42 <= _T_9260_3;
              end else begin
                if (_T_13281) begin
                  _T_16959_42 <= _T_9260_4;
                end else begin
                  if (_T_13279) begin
                    _T_16959_42 <= _T_9260_5;
                  end else begin
                    if (_T_13277) begin
                      _T_16959_42 <= _T_9260_6;
                    end else begin
                      if (_T_13275) begin
                        _T_16959_42 <= _T_9260_7;
                      end else begin
                        if (_T_13273) begin
                          _T_16959_42 <= _T_9260_8;
                        end else begin
                          if (_T_13271) begin
                            _T_16959_42 <= _T_9260_9;
                          end else begin
                            if (_T_13269) begin
                              _T_16959_42 <= _T_9260_10;
                            end else begin
                              if (_T_13267) begin
                                _T_16959_42 <= _T_9260_11;
                              end else begin
                                if (_T_13265) begin
                                  _T_16959_42 <= _T_9260_12;
                                end else begin
                                  if (_T_13263) begin
                                    _T_16959_42 <= _T_9260_13;
                                  end else begin
                                    if (_T_13261) begin
                                      _T_16959_42 <= _T_9260_14;
                                    end else begin
                                      if (_T_13259) begin
                                        _T_16959_42 <= _T_9260_15;
                                      end else begin
                                        if (_T_13257) begin
                                          _T_16959_42 <= _T_9260_16;
                                        end else begin
                                          if (_T_13255) begin
                                            _T_16959_42 <= _T_9260_17;
                                          end else begin
                                            if (_T_13253) begin
                                              _T_16959_42 <= _T_9260_18;
                                            end else begin
                                              if (_T_13251) begin
                                                _T_16959_42 <= _T_9260_19;
                                              end else begin
                                                if (_T_13249) begin
                                                  _T_16959_42 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13247) begin
                                                    _T_16959_42 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13245) begin
                                                      _T_16959_42 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13243) begin
                                                        _T_16959_42 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13241) begin
                                                          _T_16959_42 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13239) begin
                                                            _T_16959_42 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13237) begin
                                                              _T_16959_42 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13235) begin
                                                                _T_16959_42 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13233) begin
                                                                  _T_16959_42 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13231) begin
                                                                    _T_16959_42 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13229) begin
                                                                      _T_16959_42 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13227) begin
                                                                        _T_16959_42 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13225) begin
                                                                          _T_16959_42 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13223) begin
                                                                            _T_16959_42 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13221) begin
                                                                              _T_16959_42 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13219) begin
                                                                                _T_16959_42 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13217) begin
                                                                                  _T_16959_42 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13215) begin
                                                                                    _T_16959_42 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13213) begin
                                                                                      _T_16959_42 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13211) begin
                                                                                        _T_16959_42 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13209) begin
                                                                                          _T_16959_42 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13207) begin
                                                                                            _T_16959_42 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_13205) begin
                                                                                              _T_16959_42 <= _T_9260_42;
                                                                                            end else begin
                                                                                              _T_16959_42 <= 8'h0;
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_42 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_43) begin
        if (_T_13422) begin
          _T_16959_43 <= _T_9260_0;
        end else begin
          if (_T_13420) begin
            _T_16959_43 <= _T_9260_1;
          end else begin
            if (_T_13418) begin
              _T_16959_43 <= _T_9260_2;
            end else begin
              if (_T_13416) begin
                _T_16959_43 <= _T_9260_3;
              end else begin
                if (_T_13414) begin
                  _T_16959_43 <= _T_9260_4;
                end else begin
                  if (_T_13412) begin
                    _T_16959_43 <= _T_9260_5;
                  end else begin
                    if (_T_13410) begin
                      _T_16959_43 <= _T_9260_6;
                    end else begin
                      if (_T_13408) begin
                        _T_16959_43 <= _T_9260_7;
                      end else begin
                        if (_T_13406) begin
                          _T_16959_43 <= _T_9260_8;
                        end else begin
                          if (_T_13404) begin
                            _T_16959_43 <= _T_9260_9;
                          end else begin
                            if (_T_13402) begin
                              _T_16959_43 <= _T_9260_10;
                            end else begin
                              if (_T_13400) begin
                                _T_16959_43 <= _T_9260_11;
                              end else begin
                                if (_T_13398) begin
                                  _T_16959_43 <= _T_9260_12;
                                end else begin
                                  if (_T_13396) begin
                                    _T_16959_43 <= _T_9260_13;
                                  end else begin
                                    if (_T_13394) begin
                                      _T_16959_43 <= _T_9260_14;
                                    end else begin
                                      if (_T_13392) begin
                                        _T_16959_43 <= _T_9260_15;
                                      end else begin
                                        if (_T_13390) begin
                                          _T_16959_43 <= _T_9260_16;
                                        end else begin
                                          if (_T_13388) begin
                                            _T_16959_43 <= _T_9260_17;
                                          end else begin
                                            if (_T_13386) begin
                                              _T_16959_43 <= _T_9260_18;
                                            end else begin
                                              if (_T_13384) begin
                                                _T_16959_43 <= _T_9260_19;
                                              end else begin
                                                if (_T_13382) begin
                                                  _T_16959_43 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13380) begin
                                                    _T_16959_43 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13378) begin
                                                      _T_16959_43 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13376) begin
                                                        _T_16959_43 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13374) begin
                                                          _T_16959_43 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13372) begin
                                                            _T_16959_43 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13370) begin
                                                              _T_16959_43 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13368) begin
                                                                _T_16959_43 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13366) begin
                                                                  _T_16959_43 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13364) begin
                                                                    _T_16959_43 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13362) begin
                                                                      _T_16959_43 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13360) begin
                                                                        _T_16959_43 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13358) begin
                                                                          _T_16959_43 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13356) begin
                                                                            _T_16959_43 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13354) begin
                                                                              _T_16959_43 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13352) begin
                                                                                _T_16959_43 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13350) begin
                                                                                  _T_16959_43 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13348) begin
                                                                                    _T_16959_43 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13346) begin
                                                                                      _T_16959_43 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13344) begin
                                                                                        _T_16959_43 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13342) begin
                                                                                          _T_16959_43 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13340) begin
                                                                                            _T_16959_43 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_13338) begin
                                                                                              _T_16959_43 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_13336) begin
                                                                                                _T_16959_43 <= _T_9260_43;
                                                                                              end else begin
                                                                                                _T_16959_43 <= 8'h0;
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_43 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_44) begin
        if (_T_13558) begin
          _T_16959_44 <= _T_9260_0;
        end else begin
          if (_T_13556) begin
            _T_16959_44 <= _T_9260_1;
          end else begin
            if (_T_13554) begin
              _T_16959_44 <= _T_9260_2;
            end else begin
              if (_T_13552) begin
                _T_16959_44 <= _T_9260_3;
              end else begin
                if (_T_13550) begin
                  _T_16959_44 <= _T_9260_4;
                end else begin
                  if (_T_13548) begin
                    _T_16959_44 <= _T_9260_5;
                  end else begin
                    if (_T_13546) begin
                      _T_16959_44 <= _T_9260_6;
                    end else begin
                      if (_T_13544) begin
                        _T_16959_44 <= _T_9260_7;
                      end else begin
                        if (_T_13542) begin
                          _T_16959_44 <= _T_9260_8;
                        end else begin
                          if (_T_13540) begin
                            _T_16959_44 <= _T_9260_9;
                          end else begin
                            if (_T_13538) begin
                              _T_16959_44 <= _T_9260_10;
                            end else begin
                              if (_T_13536) begin
                                _T_16959_44 <= _T_9260_11;
                              end else begin
                                if (_T_13534) begin
                                  _T_16959_44 <= _T_9260_12;
                                end else begin
                                  if (_T_13532) begin
                                    _T_16959_44 <= _T_9260_13;
                                  end else begin
                                    if (_T_13530) begin
                                      _T_16959_44 <= _T_9260_14;
                                    end else begin
                                      if (_T_13528) begin
                                        _T_16959_44 <= _T_9260_15;
                                      end else begin
                                        if (_T_13526) begin
                                          _T_16959_44 <= _T_9260_16;
                                        end else begin
                                          if (_T_13524) begin
                                            _T_16959_44 <= _T_9260_17;
                                          end else begin
                                            if (_T_13522) begin
                                              _T_16959_44 <= _T_9260_18;
                                            end else begin
                                              if (_T_13520) begin
                                                _T_16959_44 <= _T_9260_19;
                                              end else begin
                                                if (_T_13518) begin
                                                  _T_16959_44 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13516) begin
                                                    _T_16959_44 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13514) begin
                                                      _T_16959_44 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13512) begin
                                                        _T_16959_44 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13510) begin
                                                          _T_16959_44 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13508) begin
                                                            _T_16959_44 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13506) begin
                                                              _T_16959_44 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13504) begin
                                                                _T_16959_44 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13502) begin
                                                                  _T_16959_44 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13500) begin
                                                                    _T_16959_44 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13498) begin
                                                                      _T_16959_44 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13496) begin
                                                                        _T_16959_44 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13494) begin
                                                                          _T_16959_44 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13492) begin
                                                                            _T_16959_44 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13490) begin
                                                                              _T_16959_44 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13488) begin
                                                                                _T_16959_44 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13486) begin
                                                                                  _T_16959_44 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13484) begin
                                                                                    _T_16959_44 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13482) begin
                                                                                      _T_16959_44 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13480) begin
                                                                                        _T_16959_44 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13478) begin
                                                                                          _T_16959_44 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13476) begin
                                                                                            _T_16959_44 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_13474) begin
                                                                                              _T_16959_44 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_13472) begin
                                                                                                _T_16959_44 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_13470) begin
                                                                                                  _T_16959_44 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  _T_16959_44 <= 8'h0;
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_44 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_45) begin
        if (_T_13697) begin
          _T_16959_45 <= _T_9260_0;
        end else begin
          if (_T_13695) begin
            _T_16959_45 <= _T_9260_1;
          end else begin
            if (_T_13693) begin
              _T_16959_45 <= _T_9260_2;
            end else begin
              if (_T_13691) begin
                _T_16959_45 <= _T_9260_3;
              end else begin
                if (_T_13689) begin
                  _T_16959_45 <= _T_9260_4;
                end else begin
                  if (_T_13687) begin
                    _T_16959_45 <= _T_9260_5;
                  end else begin
                    if (_T_13685) begin
                      _T_16959_45 <= _T_9260_6;
                    end else begin
                      if (_T_13683) begin
                        _T_16959_45 <= _T_9260_7;
                      end else begin
                        if (_T_13681) begin
                          _T_16959_45 <= _T_9260_8;
                        end else begin
                          if (_T_13679) begin
                            _T_16959_45 <= _T_9260_9;
                          end else begin
                            if (_T_13677) begin
                              _T_16959_45 <= _T_9260_10;
                            end else begin
                              if (_T_13675) begin
                                _T_16959_45 <= _T_9260_11;
                              end else begin
                                if (_T_13673) begin
                                  _T_16959_45 <= _T_9260_12;
                                end else begin
                                  if (_T_13671) begin
                                    _T_16959_45 <= _T_9260_13;
                                  end else begin
                                    if (_T_13669) begin
                                      _T_16959_45 <= _T_9260_14;
                                    end else begin
                                      if (_T_13667) begin
                                        _T_16959_45 <= _T_9260_15;
                                      end else begin
                                        if (_T_13665) begin
                                          _T_16959_45 <= _T_9260_16;
                                        end else begin
                                          if (_T_13663) begin
                                            _T_16959_45 <= _T_9260_17;
                                          end else begin
                                            if (_T_13661) begin
                                              _T_16959_45 <= _T_9260_18;
                                            end else begin
                                              if (_T_13659) begin
                                                _T_16959_45 <= _T_9260_19;
                                              end else begin
                                                if (_T_13657) begin
                                                  _T_16959_45 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13655) begin
                                                    _T_16959_45 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13653) begin
                                                      _T_16959_45 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13651) begin
                                                        _T_16959_45 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13649) begin
                                                          _T_16959_45 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13647) begin
                                                            _T_16959_45 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13645) begin
                                                              _T_16959_45 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13643) begin
                                                                _T_16959_45 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13641) begin
                                                                  _T_16959_45 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13639) begin
                                                                    _T_16959_45 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13637) begin
                                                                      _T_16959_45 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13635) begin
                                                                        _T_16959_45 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13633) begin
                                                                          _T_16959_45 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13631) begin
                                                                            _T_16959_45 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13629) begin
                                                                              _T_16959_45 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13627) begin
                                                                                _T_16959_45 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13625) begin
                                                                                  _T_16959_45 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13623) begin
                                                                                    _T_16959_45 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13621) begin
                                                                                      _T_16959_45 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13619) begin
                                                                                        _T_16959_45 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13617) begin
                                                                                          _T_16959_45 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13615) begin
                                                                                            _T_16959_45 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_13613) begin
                                                                                              _T_16959_45 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_13611) begin
                                                                                                _T_16959_45 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_13609) begin
                                                                                                  _T_16959_45 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_13607) begin
                                                                                                    _T_16959_45 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    _T_16959_45 <= 8'h0;
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_45 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_46) begin
        if (_T_13839) begin
          _T_16959_46 <= _T_9260_0;
        end else begin
          if (_T_13837) begin
            _T_16959_46 <= _T_9260_1;
          end else begin
            if (_T_13835) begin
              _T_16959_46 <= _T_9260_2;
            end else begin
              if (_T_13833) begin
                _T_16959_46 <= _T_9260_3;
              end else begin
                if (_T_13831) begin
                  _T_16959_46 <= _T_9260_4;
                end else begin
                  if (_T_13829) begin
                    _T_16959_46 <= _T_9260_5;
                  end else begin
                    if (_T_13827) begin
                      _T_16959_46 <= _T_9260_6;
                    end else begin
                      if (_T_13825) begin
                        _T_16959_46 <= _T_9260_7;
                      end else begin
                        if (_T_13823) begin
                          _T_16959_46 <= _T_9260_8;
                        end else begin
                          if (_T_13821) begin
                            _T_16959_46 <= _T_9260_9;
                          end else begin
                            if (_T_13819) begin
                              _T_16959_46 <= _T_9260_10;
                            end else begin
                              if (_T_13817) begin
                                _T_16959_46 <= _T_9260_11;
                              end else begin
                                if (_T_13815) begin
                                  _T_16959_46 <= _T_9260_12;
                                end else begin
                                  if (_T_13813) begin
                                    _T_16959_46 <= _T_9260_13;
                                  end else begin
                                    if (_T_13811) begin
                                      _T_16959_46 <= _T_9260_14;
                                    end else begin
                                      if (_T_13809) begin
                                        _T_16959_46 <= _T_9260_15;
                                      end else begin
                                        if (_T_13807) begin
                                          _T_16959_46 <= _T_9260_16;
                                        end else begin
                                          if (_T_13805) begin
                                            _T_16959_46 <= _T_9260_17;
                                          end else begin
                                            if (_T_13803) begin
                                              _T_16959_46 <= _T_9260_18;
                                            end else begin
                                              if (_T_13801) begin
                                                _T_16959_46 <= _T_9260_19;
                                              end else begin
                                                if (_T_13799) begin
                                                  _T_16959_46 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13797) begin
                                                    _T_16959_46 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13795) begin
                                                      _T_16959_46 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13793) begin
                                                        _T_16959_46 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13791) begin
                                                          _T_16959_46 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13789) begin
                                                            _T_16959_46 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13787) begin
                                                              _T_16959_46 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13785) begin
                                                                _T_16959_46 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13783) begin
                                                                  _T_16959_46 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13781) begin
                                                                    _T_16959_46 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13779) begin
                                                                      _T_16959_46 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13777) begin
                                                                        _T_16959_46 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13775) begin
                                                                          _T_16959_46 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13773) begin
                                                                            _T_16959_46 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13771) begin
                                                                              _T_16959_46 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13769) begin
                                                                                _T_16959_46 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13767) begin
                                                                                  _T_16959_46 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13765) begin
                                                                                    _T_16959_46 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13763) begin
                                                                                      _T_16959_46 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13761) begin
                                                                                        _T_16959_46 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13759) begin
                                                                                          _T_16959_46 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13757) begin
                                                                                            _T_16959_46 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_13755) begin
                                                                                              _T_16959_46 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_13753) begin
                                                                                                _T_16959_46 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_13751) begin
                                                                                                  _T_16959_46 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_13749) begin
                                                                                                    _T_16959_46 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_13747) begin
                                                                                                      _T_16959_46 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      _T_16959_46 <= 8'h0;
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_46 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_47) begin
        if (_T_13984) begin
          _T_16959_47 <= _T_9260_0;
        end else begin
          if (_T_13982) begin
            _T_16959_47 <= _T_9260_1;
          end else begin
            if (_T_13980) begin
              _T_16959_47 <= _T_9260_2;
            end else begin
              if (_T_13978) begin
                _T_16959_47 <= _T_9260_3;
              end else begin
                if (_T_13976) begin
                  _T_16959_47 <= _T_9260_4;
                end else begin
                  if (_T_13974) begin
                    _T_16959_47 <= _T_9260_5;
                  end else begin
                    if (_T_13972) begin
                      _T_16959_47 <= _T_9260_6;
                    end else begin
                      if (_T_13970) begin
                        _T_16959_47 <= _T_9260_7;
                      end else begin
                        if (_T_13968) begin
                          _T_16959_47 <= _T_9260_8;
                        end else begin
                          if (_T_13966) begin
                            _T_16959_47 <= _T_9260_9;
                          end else begin
                            if (_T_13964) begin
                              _T_16959_47 <= _T_9260_10;
                            end else begin
                              if (_T_13962) begin
                                _T_16959_47 <= _T_9260_11;
                              end else begin
                                if (_T_13960) begin
                                  _T_16959_47 <= _T_9260_12;
                                end else begin
                                  if (_T_13958) begin
                                    _T_16959_47 <= _T_9260_13;
                                  end else begin
                                    if (_T_13956) begin
                                      _T_16959_47 <= _T_9260_14;
                                    end else begin
                                      if (_T_13954) begin
                                        _T_16959_47 <= _T_9260_15;
                                      end else begin
                                        if (_T_13952) begin
                                          _T_16959_47 <= _T_9260_16;
                                        end else begin
                                          if (_T_13950) begin
                                            _T_16959_47 <= _T_9260_17;
                                          end else begin
                                            if (_T_13948) begin
                                              _T_16959_47 <= _T_9260_18;
                                            end else begin
                                              if (_T_13946) begin
                                                _T_16959_47 <= _T_9260_19;
                                              end else begin
                                                if (_T_13944) begin
                                                  _T_16959_47 <= _T_9260_20;
                                                end else begin
                                                  if (_T_13942) begin
                                                    _T_16959_47 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_13940) begin
                                                      _T_16959_47 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_13938) begin
                                                        _T_16959_47 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_13936) begin
                                                          _T_16959_47 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_13934) begin
                                                            _T_16959_47 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_13932) begin
                                                              _T_16959_47 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_13930) begin
                                                                _T_16959_47 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_13928) begin
                                                                  _T_16959_47 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_13926) begin
                                                                    _T_16959_47 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_13924) begin
                                                                      _T_16959_47 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_13922) begin
                                                                        _T_16959_47 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_13920) begin
                                                                          _T_16959_47 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_13918) begin
                                                                            _T_16959_47 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_13916) begin
                                                                              _T_16959_47 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_13914) begin
                                                                                _T_16959_47 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_13912) begin
                                                                                  _T_16959_47 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_13910) begin
                                                                                    _T_16959_47 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_13908) begin
                                                                                      _T_16959_47 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_13906) begin
                                                                                        _T_16959_47 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_13904) begin
                                                                                          _T_16959_47 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_13902) begin
                                                                                            _T_16959_47 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_13900) begin
                                                                                              _T_16959_47 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_13898) begin
                                                                                                _T_16959_47 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_13896) begin
                                                                                                  _T_16959_47 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_13894) begin
                                                                                                    _T_16959_47 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_13892) begin
                                                                                                      _T_16959_47 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_13890) begin
                                                                                                        _T_16959_47 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        _T_16959_47 <= 8'h0;
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_47 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_48) begin
        if (_T_14132) begin
          _T_16959_48 <= _T_9260_0;
        end else begin
          if (_T_14130) begin
            _T_16959_48 <= _T_9260_1;
          end else begin
            if (_T_14128) begin
              _T_16959_48 <= _T_9260_2;
            end else begin
              if (_T_14126) begin
                _T_16959_48 <= _T_9260_3;
              end else begin
                if (_T_14124) begin
                  _T_16959_48 <= _T_9260_4;
                end else begin
                  if (_T_14122) begin
                    _T_16959_48 <= _T_9260_5;
                  end else begin
                    if (_T_14120) begin
                      _T_16959_48 <= _T_9260_6;
                    end else begin
                      if (_T_14118) begin
                        _T_16959_48 <= _T_9260_7;
                      end else begin
                        if (_T_14116) begin
                          _T_16959_48 <= _T_9260_8;
                        end else begin
                          if (_T_14114) begin
                            _T_16959_48 <= _T_9260_9;
                          end else begin
                            if (_T_14112) begin
                              _T_16959_48 <= _T_9260_10;
                            end else begin
                              if (_T_14110) begin
                                _T_16959_48 <= _T_9260_11;
                              end else begin
                                if (_T_14108) begin
                                  _T_16959_48 <= _T_9260_12;
                                end else begin
                                  if (_T_14106) begin
                                    _T_16959_48 <= _T_9260_13;
                                  end else begin
                                    if (_T_14104) begin
                                      _T_16959_48 <= _T_9260_14;
                                    end else begin
                                      if (_T_14102) begin
                                        _T_16959_48 <= _T_9260_15;
                                      end else begin
                                        if (_T_14100) begin
                                          _T_16959_48 <= _T_9260_16;
                                        end else begin
                                          if (_T_14098) begin
                                            _T_16959_48 <= _T_9260_17;
                                          end else begin
                                            if (_T_14096) begin
                                              _T_16959_48 <= _T_9260_18;
                                            end else begin
                                              if (_T_14094) begin
                                                _T_16959_48 <= _T_9260_19;
                                              end else begin
                                                if (_T_14092) begin
                                                  _T_16959_48 <= _T_9260_20;
                                                end else begin
                                                  if (_T_14090) begin
                                                    _T_16959_48 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_14088) begin
                                                      _T_16959_48 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_14086) begin
                                                        _T_16959_48 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_14084) begin
                                                          _T_16959_48 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_14082) begin
                                                            _T_16959_48 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_14080) begin
                                                              _T_16959_48 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_14078) begin
                                                                _T_16959_48 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_14076) begin
                                                                  _T_16959_48 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_14074) begin
                                                                    _T_16959_48 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_14072) begin
                                                                      _T_16959_48 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_14070) begin
                                                                        _T_16959_48 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_14068) begin
                                                                          _T_16959_48 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_14066) begin
                                                                            _T_16959_48 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_14064) begin
                                                                              _T_16959_48 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_14062) begin
                                                                                _T_16959_48 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_14060) begin
                                                                                  _T_16959_48 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_14058) begin
                                                                                    _T_16959_48 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_14056) begin
                                                                                      _T_16959_48 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_14054) begin
                                                                                        _T_16959_48 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_14052) begin
                                                                                          _T_16959_48 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_14050) begin
                                                                                            _T_16959_48 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14048) begin
                                                                                              _T_16959_48 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14046) begin
                                                                                                _T_16959_48 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14044) begin
                                                                                                  _T_16959_48 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14042) begin
                                                                                                    _T_16959_48 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14040) begin
                                                                                                      _T_16959_48 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14038) begin
                                                                                                        _T_16959_48 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14036) begin
                                                                                                          _T_16959_48 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          _T_16959_48 <= 8'h0;
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_48 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_49) begin
        if (_T_14283) begin
          _T_16959_49 <= _T_9260_0;
        end else begin
          if (_T_14281) begin
            _T_16959_49 <= _T_9260_1;
          end else begin
            if (_T_14279) begin
              _T_16959_49 <= _T_9260_2;
            end else begin
              if (_T_14277) begin
                _T_16959_49 <= _T_9260_3;
              end else begin
                if (_T_14275) begin
                  _T_16959_49 <= _T_9260_4;
                end else begin
                  if (_T_14273) begin
                    _T_16959_49 <= _T_9260_5;
                  end else begin
                    if (_T_14271) begin
                      _T_16959_49 <= _T_9260_6;
                    end else begin
                      if (_T_14269) begin
                        _T_16959_49 <= _T_9260_7;
                      end else begin
                        if (_T_14267) begin
                          _T_16959_49 <= _T_9260_8;
                        end else begin
                          if (_T_14265) begin
                            _T_16959_49 <= _T_9260_9;
                          end else begin
                            if (_T_14263) begin
                              _T_16959_49 <= _T_9260_10;
                            end else begin
                              if (_T_14261) begin
                                _T_16959_49 <= _T_9260_11;
                              end else begin
                                if (_T_14259) begin
                                  _T_16959_49 <= _T_9260_12;
                                end else begin
                                  if (_T_14257) begin
                                    _T_16959_49 <= _T_9260_13;
                                  end else begin
                                    if (_T_14255) begin
                                      _T_16959_49 <= _T_9260_14;
                                    end else begin
                                      if (_T_14253) begin
                                        _T_16959_49 <= _T_9260_15;
                                      end else begin
                                        if (_T_14251) begin
                                          _T_16959_49 <= _T_9260_16;
                                        end else begin
                                          if (_T_14249) begin
                                            _T_16959_49 <= _T_9260_17;
                                          end else begin
                                            if (_T_14247) begin
                                              _T_16959_49 <= _T_9260_18;
                                            end else begin
                                              if (_T_14245) begin
                                                _T_16959_49 <= _T_9260_19;
                                              end else begin
                                                if (_T_14243) begin
                                                  _T_16959_49 <= _T_9260_20;
                                                end else begin
                                                  if (_T_14241) begin
                                                    _T_16959_49 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_14239) begin
                                                      _T_16959_49 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_14237) begin
                                                        _T_16959_49 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_14235) begin
                                                          _T_16959_49 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_14233) begin
                                                            _T_16959_49 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_14231) begin
                                                              _T_16959_49 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_14229) begin
                                                                _T_16959_49 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_14227) begin
                                                                  _T_16959_49 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_14225) begin
                                                                    _T_16959_49 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_14223) begin
                                                                      _T_16959_49 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_14221) begin
                                                                        _T_16959_49 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_14219) begin
                                                                          _T_16959_49 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_14217) begin
                                                                            _T_16959_49 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_14215) begin
                                                                              _T_16959_49 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_14213) begin
                                                                                _T_16959_49 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_14211) begin
                                                                                  _T_16959_49 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_14209) begin
                                                                                    _T_16959_49 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_14207) begin
                                                                                      _T_16959_49 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_14205) begin
                                                                                        _T_16959_49 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_14203) begin
                                                                                          _T_16959_49 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_14201) begin
                                                                                            _T_16959_49 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14199) begin
                                                                                              _T_16959_49 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14197) begin
                                                                                                _T_16959_49 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14195) begin
                                                                                                  _T_16959_49 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14193) begin
                                                                                                    _T_16959_49 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14191) begin
                                                                                                      _T_16959_49 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14189) begin
                                                                                                        _T_16959_49 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14187) begin
                                                                                                          _T_16959_49 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_14185) begin
                                                                                                            _T_16959_49 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            _T_16959_49 <= 8'h0;
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_49 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_50) begin
        if (_T_14437) begin
          _T_16959_50 <= _T_9260_0;
        end else begin
          if (_T_14435) begin
            _T_16959_50 <= _T_9260_1;
          end else begin
            if (_T_14433) begin
              _T_16959_50 <= _T_9260_2;
            end else begin
              if (_T_14431) begin
                _T_16959_50 <= _T_9260_3;
              end else begin
                if (_T_14429) begin
                  _T_16959_50 <= _T_9260_4;
                end else begin
                  if (_T_14427) begin
                    _T_16959_50 <= _T_9260_5;
                  end else begin
                    if (_T_14425) begin
                      _T_16959_50 <= _T_9260_6;
                    end else begin
                      if (_T_14423) begin
                        _T_16959_50 <= _T_9260_7;
                      end else begin
                        if (_T_14421) begin
                          _T_16959_50 <= _T_9260_8;
                        end else begin
                          if (_T_14419) begin
                            _T_16959_50 <= _T_9260_9;
                          end else begin
                            if (_T_14417) begin
                              _T_16959_50 <= _T_9260_10;
                            end else begin
                              if (_T_14415) begin
                                _T_16959_50 <= _T_9260_11;
                              end else begin
                                if (_T_14413) begin
                                  _T_16959_50 <= _T_9260_12;
                                end else begin
                                  if (_T_14411) begin
                                    _T_16959_50 <= _T_9260_13;
                                  end else begin
                                    if (_T_14409) begin
                                      _T_16959_50 <= _T_9260_14;
                                    end else begin
                                      if (_T_14407) begin
                                        _T_16959_50 <= _T_9260_15;
                                      end else begin
                                        if (_T_14405) begin
                                          _T_16959_50 <= _T_9260_16;
                                        end else begin
                                          if (_T_14403) begin
                                            _T_16959_50 <= _T_9260_17;
                                          end else begin
                                            if (_T_14401) begin
                                              _T_16959_50 <= _T_9260_18;
                                            end else begin
                                              if (_T_14399) begin
                                                _T_16959_50 <= _T_9260_19;
                                              end else begin
                                                if (_T_14397) begin
                                                  _T_16959_50 <= _T_9260_20;
                                                end else begin
                                                  if (_T_14395) begin
                                                    _T_16959_50 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_14393) begin
                                                      _T_16959_50 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_14391) begin
                                                        _T_16959_50 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_14389) begin
                                                          _T_16959_50 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_14387) begin
                                                            _T_16959_50 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_14385) begin
                                                              _T_16959_50 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_14383) begin
                                                                _T_16959_50 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_14381) begin
                                                                  _T_16959_50 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_14379) begin
                                                                    _T_16959_50 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_14377) begin
                                                                      _T_16959_50 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_14375) begin
                                                                        _T_16959_50 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_14373) begin
                                                                          _T_16959_50 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_14371) begin
                                                                            _T_16959_50 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_14369) begin
                                                                              _T_16959_50 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_14367) begin
                                                                                _T_16959_50 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_14365) begin
                                                                                  _T_16959_50 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_14363) begin
                                                                                    _T_16959_50 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_14361) begin
                                                                                      _T_16959_50 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_14359) begin
                                                                                        _T_16959_50 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_14357) begin
                                                                                          _T_16959_50 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_14355) begin
                                                                                            _T_16959_50 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14353) begin
                                                                                              _T_16959_50 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14351) begin
                                                                                                _T_16959_50 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14349) begin
                                                                                                  _T_16959_50 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14347) begin
                                                                                                    _T_16959_50 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14345) begin
                                                                                                      _T_16959_50 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14343) begin
                                                                                                        _T_16959_50 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14341) begin
                                                                                                          _T_16959_50 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_14339) begin
                                                                                                            _T_16959_50 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_14337) begin
                                                                                                              _T_16959_50 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              _T_16959_50 <= 8'h0;
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_50 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_51) begin
        if (_T_14594) begin
          _T_16959_51 <= _T_9260_0;
        end else begin
          if (_T_14592) begin
            _T_16959_51 <= _T_9260_1;
          end else begin
            if (_T_14590) begin
              _T_16959_51 <= _T_9260_2;
            end else begin
              if (_T_14588) begin
                _T_16959_51 <= _T_9260_3;
              end else begin
                if (_T_14586) begin
                  _T_16959_51 <= _T_9260_4;
                end else begin
                  if (_T_14584) begin
                    _T_16959_51 <= _T_9260_5;
                  end else begin
                    if (_T_14582) begin
                      _T_16959_51 <= _T_9260_6;
                    end else begin
                      if (_T_14580) begin
                        _T_16959_51 <= _T_9260_7;
                      end else begin
                        if (_T_14578) begin
                          _T_16959_51 <= _T_9260_8;
                        end else begin
                          if (_T_14576) begin
                            _T_16959_51 <= _T_9260_9;
                          end else begin
                            if (_T_14574) begin
                              _T_16959_51 <= _T_9260_10;
                            end else begin
                              if (_T_14572) begin
                                _T_16959_51 <= _T_9260_11;
                              end else begin
                                if (_T_14570) begin
                                  _T_16959_51 <= _T_9260_12;
                                end else begin
                                  if (_T_14568) begin
                                    _T_16959_51 <= _T_9260_13;
                                  end else begin
                                    if (_T_14566) begin
                                      _T_16959_51 <= _T_9260_14;
                                    end else begin
                                      if (_T_14564) begin
                                        _T_16959_51 <= _T_9260_15;
                                      end else begin
                                        if (_T_14562) begin
                                          _T_16959_51 <= _T_9260_16;
                                        end else begin
                                          if (_T_14560) begin
                                            _T_16959_51 <= _T_9260_17;
                                          end else begin
                                            if (_T_14558) begin
                                              _T_16959_51 <= _T_9260_18;
                                            end else begin
                                              if (_T_14556) begin
                                                _T_16959_51 <= _T_9260_19;
                                              end else begin
                                                if (_T_14554) begin
                                                  _T_16959_51 <= _T_9260_20;
                                                end else begin
                                                  if (_T_14552) begin
                                                    _T_16959_51 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_14550) begin
                                                      _T_16959_51 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_14548) begin
                                                        _T_16959_51 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_14546) begin
                                                          _T_16959_51 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_14544) begin
                                                            _T_16959_51 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_14542) begin
                                                              _T_16959_51 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_14540) begin
                                                                _T_16959_51 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_14538) begin
                                                                  _T_16959_51 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_14536) begin
                                                                    _T_16959_51 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_14534) begin
                                                                      _T_16959_51 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_14532) begin
                                                                        _T_16959_51 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_14530) begin
                                                                          _T_16959_51 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_14528) begin
                                                                            _T_16959_51 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_14526) begin
                                                                              _T_16959_51 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_14524) begin
                                                                                _T_16959_51 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_14522) begin
                                                                                  _T_16959_51 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_14520) begin
                                                                                    _T_16959_51 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_14518) begin
                                                                                      _T_16959_51 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_14516) begin
                                                                                        _T_16959_51 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_14514) begin
                                                                                          _T_16959_51 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_14512) begin
                                                                                            _T_16959_51 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14510) begin
                                                                                              _T_16959_51 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14508) begin
                                                                                                _T_16959_51 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14506) begin
                                                                                                  _T_16959_51 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14504) begin
                                                                                                    _T_16959_51 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14502) begin
                                                                                                      _T_16959_51 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14500) begin
                                                                                                        _T_16959_51 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14498) begin
                                                                                                          _T_16959_51 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_14496) begin
                                                                                                            _T_16959_51 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_14494) begin
                                                                                                              _T_16959_51 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_14492) begin
                                                                                                                _T_16959_51 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                _T_16959_51 <= 8'h0;
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_51 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_52) begin
        if (_T_14754) begin
          _T_16959_52 <= _T_9260_0;
        end else begin
          if (_T_14752) begin
            _T_16959_52 <= _T_9260_1;
          end else begin
            if (_T_14750) begin
              _T_16959_52 <= _T_9260_2;
            end else begin
              if (_T_14748) begin
                _T_16959_52 <= _T_9260_3;
              end else begin
                if (_T_14746) begin
                  _T_16959_52 <= _T_9260_4;
                end else begin
                  if (_T_14744) begin
                    _T_16959_52 <= _T_9260_5;
                  end else begin
                    if (_T_14742) begin
                      _T_16959_52 <= _T_9260_6;
                    end else begin
                      if (_T_14740) begin
                        _T_16959_52 <= _T_9260_7;
                      end else begin
                        if (_T_14738) begin
                          _T_16959_52 <= _T_9260_8;
                        end else begin
                          if (_T_14736) begin
                            _T_16959_52 <= _T_9260_9;
                          end else begin
                            if (_T_14734) begin
                              _T_16959_52 <= _T_9260_10;
                            end else begin
                              if (_T_14732) begin
                                _T_16959_52 <= _T_9260_11;
                              end else begin
                                if (_T_14730) begin
                                  _T_16959_52 <= _T_9260_12;
                                end else begin
                                  if (_T_14728) begin
                                    _T_16959_52 <= _T_9260_13;
                                  end else begin
                                    if (_T_14726) begin
                                      _T_16959_52 <= _T_9260_14;
                                    end else begin
                                      if (_T_14724) begin
                                        _T_16959_52 <= _T_9260_15;
                                      end else begin
                                        if (_T_14722) begin
                                          _T_16959_52 <= _T_9260_16;
                                        end else begin
                                          if (_T_14720) begin
                                            _T_16959_52 <= _T_9260_17;
                                          end else begin
                                            if (_T_14718) begin
                                              _T_16959_52 <= _T_9260_18;
                                            end else begin
                                              if (_T_14716) begin
                                                _T_16959_52 <= _T_9260_19;
                                              end else begin
                                                if (_T_14714) begin
                                                  _T_16959_52 <= _T_9260_20;
                                                end else begin
                                                  if (_T_14712) begin
                                                    _T_16959_52 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_14710) begin
                                                      _T_16959_52 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_14708) begin
                                                        _T_16959_52 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_14706) begin
                                                          _T_16959_52 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_14704) begin
                                                            _T_16959_52 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_14702) begin
                                                              _T_16959_52 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_14700) begin
                                                                _T_16959_52 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_14698) begin
                                                                  _T_16959_52 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_14696) begin
                                                                    _T_16959_52 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_14694) begin
                                                                      _T_16959_52 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_14692) begin
                                                                        _T_16959_52 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_14690) begin
                                                                          _T_16959_52 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_14688) begin
                                                                            _T_16959_52 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_14686) begin
                                                                              _T_16959_52 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_14684) begin
                                                                                _T_16959_52 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_14682) begin
                                                                                  _T_16959_52 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_14680) begin
                                                                                    _T_16959_52 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_14678) begin
                                                                                      _T_16959_52 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_14676) begin
                                                                                        _T_16959_52 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_14674) begin
                                                                                          _T_16959_52 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_14672) begin
                                                                                            _T_16959_52 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14670) begin
                                                                                              _T_16959_52 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14668) begin
                                                                                                _T_16959_52 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14666) begin
                                                                                                  _T_16959_52 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14664) begin
                                                                                                    _T_16959_52 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14662) begin
                                                                                                      _T_16959_52 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14660) begin
                                                                                                        _T_16959_52 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14658) begin
                                                                                                          _T_16959_52 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_14656) begin
                                                                                                            _T_16959_52 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_14654) begin
                                                                                                              _T_16959_52 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_14652) begin
                                                                                                                _T_16959_52 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_14650) begin
                                                                                                                  _T_16959_52 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  _T_16959_52 <= 8'h0;
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_52 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_53) begin
        if (_T_14917) begin
          _T_16959_53 <= _T_9260_0;
        end else begin
          if (_T_14915) begin
            _T_16959_53 <= _T_9260_1;
          end else begin
            if (_T_14913) begin
              _T_16959_53 <= _T_9260_2;
            end else begin
              if (_T_14911) begin
                _T_16959_53 <= _T_9260_3;
              end else begin
                if (_T_14909) begin
                  _T_16959_53 <= _T_9260_4;
                end else begin
                  if (_T_14907) begin
                    _T_16959_53 <= _T_9260_5;
                  end else begin
                    if (_T_14905) begin
                      _T_16959_53 <= _T_9260_6;
                    end else begin
                      if (_T_14903) begin
                        _T_16959_53 <= _T_9260_7;
                      end else begin
                        if (_T_14901) begin
                          _T_16959_53 <= _T_9260_8;
                        end else begin
                          if (_T_14899) begin
                            _T_16959_53 <= _T_9260_9;
                          end else begin
                            if (_T_14897) begin
                              _T_16959_53 <= _T_9260_10;
                            end else begin
                              if (_T_14895) begin
                                _T_16959_53 <= _T_9260_11;
                              end else begin
                                if (_T_14893) begin
                                  _T_16959_53 <= _T_9260_12;
                                end else begin
                                  if (_T_14891) begin
                                    _T_16959_53 <= _T_9260_13;
                                  end else begin
                                    if (_T_14889) begin
                                      _T_16959_53 <= _T_9260_14;
                                    end else begin
                                      if (_T_14887) begin
                                        _T_16959_53 <= _T_9260_15;
                                      end else begin
                                        if (_T_14885) begin
                                          _T_16959_53 <= _T_9260_16;
                                        end else begin
                                          if (_T_14883) begin
                                            _T_16959_53 <= _T_9260_17;
                                          end else begin
                                            if (_T_14881) begin
                                              _T_16959_53 <= _T_9260_18;
                                            end else begin
                                              if (_T_14879) begin
                                                _T_16959_53 <= _T_9260_19;
                                              end else begin
                                                if (_T_14877) begin
                                                  _T_16959_53 <= _T_9260_20;
                                                end else begin
                                                  if (_T_14875) begin
                                                    _T_16959_53 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_14873) begin
                                                      _T_16959_53 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_14871) begin
                                                        _T_16959_53 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_14869) begin
                                                          _T_16959_53 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_14867) begin
                                                            _T_16959_53 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_14865) begin
                                                              _T_16959_53 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_14863) begin
                                                                _T_16959_53 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_14861) begin
                                                                  _T_16959_53 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_14859) begin
                                                                    _T_16959_53 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_14857) begin
                                                                      _T_16959_53 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_14855) begin
                                                                        _T_16959_53 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_14853) begin
                                                                          _T_16959_53 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_14851) begin
                                                                            _T_16959_53 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_14849) begin
                                                                              _T_16959_53 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_14847) begin
                                                                                _T_16959_53 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_14845) begin
                                                                                  _T_16959_53 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_14843) begin
                                                                                    _T_16959_53 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_14841) begin
                                                                                      _T_16959_53 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_14839) begin
                                                                                        _T_16959_53 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_14837) begin
                                                                                          _T_16959_53 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_14835) begin
                                                                                            _T_16959_53 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14833) begin
                                                                                              _T_16959_53 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14831) begin
                                                                                                _T_16959_53 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14829) begin
                                                                                                  _T_16959_53 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14827) begin
                                                                                                    _T_16959_53 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14825) begin
                                                                                                      _T_16959_53 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14823) begin
                                                                                                        _T_16959_53 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14821) begin
                                                                                                          _T_16959_53 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_14819) begin
                                                                                                            _T_16959_53 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_14817) begin
                                                                                                              _T_16959_53 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_14815) begin
                                                                                                                _T_16959_53 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_14813) begin
                                                                                                                  _T_16959_53 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_14811) begin
                                                                                                                    _T_16959_53 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    _T_16959_53 <= 8'h0;
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_53 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_54) begin
        if (_T_15083) begin
          _T_16959_54 <= _T_9260_0;
        end else begin
          if (_T_15081) begin
            _T_16959_54 <= _T_9260_1;
          end else begin
            if (_T_15079) begin
              _T_16959_54 <= _T_9260_2;
            end else begin
              if (_T_15077) begin
                _T_16959_54 <= _T_9260_3;
              end else begin
                if (_T_15075) begin
                  _T_16959_54 <= _T_9260_4;
                end else begin
                  if (_T_15073) begin
                    _T_16959_54 <= _T_9260_5;
                  end else begin
                    if (_T_15071) begin
                      _T_16959_54 <= _T_9260_6;
                    end else begin
                      if (_T_15069) begin
                        _T_16959_54 <= _T_9260_7;
                      end else begin
                        if (_T_15067) begin
                          _T_16959_54 <= _T_9260_8;
                        end else begin
                          if (_T_15065) begin
                            _T_16959_54 <= _T_9260_9;
                          end else begin
                            if (_T_15063) begin
                              _T_16959_54 <= _T_9260_10;
                            end else begin
                              if (_T_15061) begin
                                _T_16959_54 <= _T_9260_11;
                              end else begin
                                if (_T_15059) begin
                                  _T_16959_54 <= _T_9260_12;
                                end else begin
                                  if (_T_15057) begin
                                    _T_16959_54 <= _T_9260_13;
                                  end else begin
                                    if (_T_15055) begin
                                      _T_16959_54 <= _T_9260_14;
                                    end else begin
                                      if (_T_15053) begin
                                        _T_16959_54 <= _T_9260_15;
                                      end else begin
                                        if (_T_15051) begin
                                          _T_16959_54 <= _T_9260_16;
                                        end else begin
                                          if (_T_15049) begin
                                            _T_16959_54 <= _T_9260_17;
                                          end else begin
                                            if (_T_15047) begin
                                              _T_16959_54 <= _T_9260_18;
                                            end else begin
                                              if (_T_15045) begin
                                                _T_16959_54 <= _T_9260_19;
                                              end else begin
                                                if (_T_15043) begin
                                                  _T_16959_54 <= _T_9260_20;
                                                end else begin
                                                  if (_T_15041) begin
                                                    _T_16959_54 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_15039) begin
                                                      _T_16959_54 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_15037) begin
                                                        _T_16959_54 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_15035) begin
                                                          _T_16959_54 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_15033) begin
                                                            _T_16959_54 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_15031) begin
                                                              _T_16959_54 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_15029) begin
                                                                _T_16959_54 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_15027) begin
                                                                  _T_16959_54 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_15025) begin
                                                                    _T_16959_54 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_15023) begin
                                                                      _T_16959_54 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_15021) begin
                                                                        _T_16959_54 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_15019) begin
                                                                          _T_16959_54 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_15017) begin
                                                                            _T_16959_54 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_15015) begin
                                                                              _T_16959_54 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_15013) begin
                                                                                _T_16959_54 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_15011) begin
                                                                                  _T_16959_54 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_15009) begin
                                                                                    _T_16959_54 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_15007) begin
                                                                                      _T_16959_54 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_15005) begin
                                                                                        _T_16959_54 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_15003) begin
                                                                                          _T_16959_54 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_15001) begin
                                                                                            _T_16959_54 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_14999) begin
                                                                                              _T_16959_54 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_14997) begin
                                                                                                _T_16959_54 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_14995) begin
                                                                                                  _T_16959_54 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_14993) begin
                                                                                                    _T_16959_54 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_14991) begin
                                                                                                      _T_16959_54 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_14989) begin
                                                                                                        _T_16959_54 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_14987) begin
                                                                                                          _T_16959_54 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_14985) begin
                                                                                                            _T_16959_54 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_14983) begin
                                                                                                              _T_16959_54 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_14981) begin
                                                                                                                _T_16959_54 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_14979) begin
                                                                                                                  _T_16959_54 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_14977) begin
                                                                                                                    _T_16959_54 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_14975) begin
                                                                                                                      _T_16959_54 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      _T_16959_54 <= 8'h0;
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_54 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_55) begin
        if (_T_15252) begin
          _T_16959_55 <= _T_9260_0;
        end else begin
          if (_T_15250) begin
            _T_16959_55 <= _T_9260_1;
          end else begin
            if (_T_15248) begin
              _T_16959_55 <= _T_9260_2;
            end else begin
              if (_T_15246) begin
                _T_16959_55 <= _T_9260_3;
              end else begin
                if (_T_15244) begin
                  _T_16959_55 <= _T_9260_4;
                end else begin
                  if (_T_15242) begin
                    _T_16959_55 <= _T_9260_5;
                  end else begin
                    if (_T_15240) begin
                      _T_16959_55 <= _T_9260_6;
                    end else begin
                      if (_T_15238) begin
                        _T_16959_55 <= _T_9260_7;
                      end else begin
                        if (_T_15236) begin
                          _T_16959_55 <= _T_9260_8;
                        end else begin
                          if (_T_15234) begin
                            _T_16959_55 <= _T_9260_9;
                          end else begin
                            if (_T_15232) begin
                              _T_16959_55 <= _T_9260_10;
                            end else begin
                              if (_T_15230) begin
                                _T_16959_55 <= _T_9260_11;
                              end else begin
                                if (_T_15228) begin
                                  _T_16959_55 <= _T_9260_12;
                                end else begin
                                  if (_T_15226) begin
                                    _T_16959_55 <= _T_9260_13;
                                  end else begin
                                    if (_T_15224) begin
                                      _T_16959_55 <= _T_9260_14;
                                    end else begin
                                      if (_T_15222) begin
                                        _T_16959_55 <= _T_9260_15;
                                      end else begin
                                        if (_T_15220) begin
                                          _T_16959_55 <= _T_9260_16;
                                        end else begin
                                          if (_T_15218) begin
                                            _T_16959_55 <= _T_9260_17;
                                          end else begin
                                            if (_T_15216) begin
                                              _T_16959_55 <= _T_9260_18;
                                            end else begin
                                              if (_T_15214) begin
                                                _T_16959_55 <= _T_9260_19;
                                              end else begin
                                                if (_T_15212) begin
                                                  _T_16959_55 <= _T_9260_20;
                                                end else begin
                                                  if (_T_15210) begin
                                                    _T_16959_55 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_15208) begin
                                                      _T_16959_55 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_15206) begin
                                                        _T_16959_55 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_15204) begin
                                                          _T_16959_55 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_15202) begin
                                                            _T_16959_55 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_15200) begin
                                                              _T_16959_55 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_15198) begin
                                                                _T_16959_55 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_15196) begin
                                                                  _T_16959_55 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_15194) begin
                                                                    _T_16959_55 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_15192) begin
                                                                      _T_16959_55 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_15190) begin
                                                                        _T_16959_55 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_15188) begin
                                                                          _T_16959_55 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_15186) begin
                                                                            _T_16959_55 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_15184) begin
                                                                              _T_16959_55 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_15182) begin
                                                                                _T_16959_55 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_15180) begin
                                                                                  _T_16959_55 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_15178) begin
                                                                                    _T_16959_55 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_15176) begin
                                                                                      _T_16959_55 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_15174) begin
                                                                                        _T_16959_55 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_15172) begin
                                                                                          _T_16959_55 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_15170) begin
                                                                                            _T_16959_55 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_15168) begin
                                                                                              _T_16959_55 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_15166) begin
                                                                                                _T_16959_55 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_15164) begin
                                                                                                  _T_16959_55 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_15162) begin
                                                                                                    _T_16959_55 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_15160) begin
                                                                                                      _T_16959_55 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_15158) begin
                                                                                                        _T_16959_55 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_15156) begin
                                                                                                          _T_16959_55 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_15154) begin
                                                                                                            _T_16959_55 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_15152) begin
                                                                                                              _T_16959_55 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_15150) begin
                                                                                                                _T_16959_55 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_15148) begin
                                                                                                                  _T_16959_55 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15146) begin
                                                                                                                    _T_16959_55 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_15144) begin
                                                                                                                      _T_16959_55 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_15142) begin
                                                                                                                        _T_16959_55 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        _T_16959_55 <= 8'h0;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_55 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_56) begin
        if (_T_15424) begin
          _T_16959_56 <= _T_9260_0;
        end else begin
          if (_T_15422) begin
            _T_16959_56 <= _T_9260_1;
          end else begin
            if (_T_15420) begin
              _T_16959_56 <= _T_9260_2;
            end else begin
              if (_T_15418) begin
                _T_16959_56 <= _T_9260_3;
              end else begin
                if (_T_15416) begin
                  _T_16959_56 <= _T_9260_4;
                end else begin
                  if (_T_15414) begin
                    _T_16959_56 <= _T_9260_5;
                  end else begin
                    if (_T_15412) begin
                      _T_16959_56 <= _T_9260_6;
                    end else begin
                      if (_T_15410) begin
                        _T_16959_56 <= _T_9260_7;
                      end else begin
                        if (_T_15408) begin
                          _T_16959_56 <= _T_9260_8;
                        end else begin
                          if (_T_15406) begin
                            _T_16959_56 <= _T_9260_9;
                          end else begin
                            if (_T_15404) begin
                              _T_16959_56 <= _T_9260_10;
                            end else begin
                              if (_T_15402) begin
                                _T_16959_56 <= _T_9260_11;
                              end else begin
                                if (_T_15400) begin
                                  _T_16959_56 <= _T_9260_12;
                                end else begin
                                  if (_T_15398) begin
                                    _T_16959_56 <= _T_9260_13;
                                  end else begin
                                    if (_T_15396) begin
                                      _T_16959_56 <= _T_9260_14;
                                    end else begin
                                      if (_T_15394) begin
                                        _T_16959_56 <= _T_9260_15;
                                      end else begin
                                        if (_T_15392) begin
                                          _T_16959_56 <= _T_9260_16;
                                        end else begin
                                          if (_T_15390) begin
                                            _T_16959_56 <= _T_9260_17;
                                          end else begin
                                            if (_T_15388) begin
                                              _T_16959_56 <= _T_9260_18;
                                            end else begin
                                              if (_T_15386) begin
                                                _T_16959_56 <= _T_9260_19;
                                              end else begin
                                                if (_T_15384) begin
                                                  _T_16959_56 <= _T_9260_20;
                                                end else begin
                                                  if (_T_15382) begin
                                                    _T_16959_56 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_15380) begin
                                                      _T_16959_56 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_15378) begin
                                                        _T_16959_56 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_15376) begin
                                                          _T_16959_56 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_15374) begin
                                                            _T_16959_56 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_15372) begin
                                                              _T_16959_56 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_15370) begin
                                                                _T_16959_56 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_15368) begin
                                                                  _T_16959_56 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_15366) begin
                                                                    _T_16959_56 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_15364) begin
                                                                      _T_16959_56 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_15362) begin
                                                                        _T_16959_56 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_15360) begin
                                                                          _T_16959_56 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_15358) begin
                                                                            _T_16959_56 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_15356) begin
                                                                              _T_16959_56 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_15354) begin
                                                                                _T_16959_56 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_15352) begin
                                                                                  _T_16959_56 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_15350) begin
                                                                                    _T_16959_56 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_15348) begin
                                                                                      _T_16959_56 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_15346) begin
                                                                                        _T_16959_56 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_15344) begin
                                                                                          _T_16959_56 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_15342) begin
                                                                                            _T_16959_56 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_15340) begin
                                                                                              _T_16959_56 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_15338) begin
                                                                                                _T_16959_56 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_15336) begin
                                                                                                  _T_16959_56 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_15334) begin
                                                                                                    _T_16959_56 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_15332) begin
                                                                                                      _T_16959_56 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_15330) begin
                                                                                                        _T_16959_56 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_15328) begin
                                                                                                          _T_16959_56 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_15326) begin
                                                                                                            _T_16959_56 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_15324) begin
                                                                                                              _T_16959_56 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_15322) begin
                                                                                                                _T_16959_56 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_15320) begin
                                                                                                                  _T_16959_56 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15318) begin
                                                                                                                    _T_16959_56 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_15316) begin
                                                                                                                      _T_16959_56 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_15314) begin
                                                                                                                        _T_16959_56 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_15312) begin
                                                                                                                          _T_16959_56 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          _T_16959_56 <= 8'h0;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_56 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_57) begin
        if (_T_15599) begin
          _T_16959_57 <= _T_9260_0;
        end else begin
          if (_T_15597) begin
            _T_16959_57 <= _T_9260_1;
          end else begin
            if (_T_15595) begin
              _T_16959_57 <= _T_9260_2;
            end else begin
              if (_T_15593) begin
                _T_16959_57 <= _T_9260_3;
              end else begin
                if (_T_15591) begin
                  _T_16959_57 <= _T_9260_4;
                end else begin
                  if (_T_15589) begin
                    _T_16959_57 <= _T_9260_5;
                  end else begin
                    if (_T_15587) begin
                      _T_16959_57 <= _T_9260_6;
                    end else begin
                      if (_T_15585) begin
                        _T_16959_57 <= _T_9260_7;
                      end else begin
                        if (_T_15583) begin
                          _T_16959_57 <= _T_9260_8;
                        end else begin
                          if (_T_15581) begin
                            _T_16959_57 <= _T_9260_9;
                          end else begin
                            if (_T_15579) begin
                              _T_16959_57 <= _T_9260_10;
                            end else begin
                              if (_T_15577) begin
                                _T_16959_57 <= _T_9260_11;
                              end else begin
                                if (_T_15575) begin
                                  _T_16959_57 <= _T_9260_12;
                                end else begin
                                  if (_T_15573) begin
                                    _T_16959_57 <= _T_9260_13;
                                  end else begin
                                    if (_T_15571) begin
                                      _T_16959_57 <= _T_9260_14;
                                    end else begin
                                      if (_T_15569) begin
                                        _T_16959_57 <= _T_9260_15;
                                      end else begin
                                        if (_T_15567) begin
                                          _T_16959_57 <= _T_9260_16;
                                        end else begin
                                          if (_T_15565) begin
                                            _T_16959_57 <= _T_9260_17;
                                          end else begin
                                            if (_T_15563) begin
                                              _T_16959_57 <= _T_9260_18;
                                            end else begin
                                              if (_T_15561) begin
                                                _T_16959_57 <= _T_9260_19;
                                              end else begin
                                                if (_T_15559) begin
                                                  _T_16959_57 <= _T_9260_20;
                                                end else begin
                                                  if (_T_15557) begin
                                                    _T_16959_57 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_15555) begin
                                                      _T_16959_57 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_15553) begin
                                                        _T_16959_57 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_15551) begin
                                                          _T_16959_57 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_15549) begin
                                                            _T_16959_57 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_15547) begin
                                                              _T_16959_57 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_15545) begin
                                                                _T_16959_57 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_15543) begin
                                                                  _T_16959_57 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_15541) begin
                                                                    _T_16959_57 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_15539) begin
                                                                      _T_16959_57 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_15537) begin
                                                                        _T_16959_57 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_15535) begin
                                                                          _T_16959_57 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_15533) begin
                                                                            _T_16959_57 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_15531) begin
                                                                              _T_16959_57 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_15529) begin
                                                                                _T_16959_57 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_15527) begin
                                                                                  _T_16959_57 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_15525) begin
                                                                                    _T_16959_57 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_15523) begin
                                                                                      _T_16959_57 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_15521) begin
                                                                                        _T_16959_57 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_15519) begin
                                                                                          _T_16959_57 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_15517) begin
                                                                                            _T_16959_57 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_15515) begin
                                                                                              _T_16959_57 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_15513) begin
                                                                                                _T_16959_57 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_15511) begin
                                                                                                  _T_16959_57 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_15509) begin
                                                                                                    _T_16959_57 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_15507) begin
                                                                                                      _T_16959_57 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_15505) begin
                                                                                                        _T_16959_57 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_15503) begin
                                                                                                          _T_16959_57 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_15501) begin
                                                                                                            _T_16959_57 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_15499) begin
                                                                                                              _T_16959_57 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_15497) begin
                                                                                                                _T_16959_57 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_15495) begin
                                                                                                                  _T_16959_57 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15493) begin
                                                                                                                    _T_16959_57 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_15491) begin
                                                                                                                      _T_16959_57 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_15489) begin
                                                                                                                        _T_16959_57 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_15487) begin
                                                                                                                          _T_16959_57 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_15485) begin
                                                                                                                            _T_16959_57 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            _T_16959_57 <= 8'h0;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_57 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_58) begin
        if (_T_15777) begin
          _T_16959_58 <= _T_9260_0;
        end else begin
          if (_T_15775) begin
            _T_16959_58 <= _T_9260_1;
          end else begin
            if (_T_15773) begin
              _T_16959_58 <= _T_9260_2;
            end else begin
              if (_T_15771) begin
                _T_16959_58 <= _T_9260_3;
              end else begin
                if (_T_15769) begin
                  _T_16959_58 <= _T_9260_4;
                end else begin
                  if (_T_15767) begin
                    _T_16959_58 <= _T_9260_5;
                  end else begin
                    if (_T_15765) begin
                      _T_16959_58 <= _T_9260_6;
                    end else begin
                      if (_T_15763) begin
                        _T_16959_58 <= _T_9260_7;
                      end else begin
                        if (_T_15761) begin
                          _T_16959_58 <= _T_9260_8;
                        end else begin
                          if (_T_15759) begin
                            _T_16959_58 <= _T_9260_9;
                          end else begin
                            if (_T_15757) begin
                              _T_16959_58 <= _T_9260_10;
                            end else begin
                              if (_T_15755) begin
                                _T_16959_58 <= _T_9260_11;
                              end else begin
                                if (_T_15753) begin
                                  _T_16959_58 <= _T_9260_12;
                                end else begin
                                  if (_T_15751) begin
                                    _T_16959_58 <= _T_9260_13;
                                  end else begin
                                    if (_T_15749) begin
                                      _T_16959_58 <= _T_9260_14;
                                    end else begin
                                      if (_T_15747) begin
                                        _T_16959_58 <= _T_9260_15;
                                      end else begin
                                        if (_T_15745) begin
                                          _T_16959_58 <= _T_9260_16;
                                        end else begin
                                          if (_T_15743) begin
                                            _T_16959_58 <= _T_9260_17;
                                          end else begin
                                            if (_T_15741) begin
                                              _T_16959_58 <= _T_9260_18;
                                            end else begin
                                              if (_T_15739) begin
                                                _T_16959_58 <= _T_9260_19;
                                              end else begin
                                                if (_T_15737) begin
                                                  _T_16959_58 <= _T_9260_20;
                                                end else begin
                                                  if (_T_15735) begin
                                                    _T_16959_58 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_15733) begin
                                                      _T_16959_58 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_15731) begin
                                                        _T_16959_58 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_15729) begin
                                                          _T_16959_58 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_15727) begin
                                                            _T_16959_58 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_15725) begin
                                                              _T_16959_58 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_15723) begin
                                                                _T_16959_58 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_15721) begin
                                                                  _T_16959_58 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_15719) begin
                                                                    _T_16959_58 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_15717) begin
                                                                      _T_16959_58 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_15715) begin
                                                                        _T_16959_58 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_15713) begin
                                                                          _T_16959_58 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_15711) begin
                                                                            _T_16959_58 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_15709) begin
                                                                              _T_16959_58 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_15707) begin
                                                                                _T_16959_58 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_15705) begin
                                                                                  _T_16959_58 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_15703) begin
                                                                                    _T_16959_58 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_15701) begin
                                                                                      _T_16959_58 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_15699) begin
                                                                                        _T_16959_58 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_15697) begin
                                                                                          _T_16959_58 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_15695) begin
                                                                                            _T_16959_58 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_15693) begin
                                                                                              _T_16959_58 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_15691) begin
                                                                                                _T_16959_58 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_15689) begin
                                                                                                  _T_16959_58 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_15687) begin
                                                                                                    _T_16959_58 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_15685) begin
                                                                                                      _T_16959_58 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_15683) begin
                                                                                                        _T_16959_58 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_15681) begin
                                                                                                          _T_16959_58 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_15679) begin
                                                                                                            _T_16959_58 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_15677) begin
                                                                                                              _T_16959_58 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_15675) begin
                                                                                                                _T_16959_58 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_15673) begin
                                                                                                                  _T_16959_58 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15671) begin
                                                                                                                    _T_16959_58 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_15669) begin
                                                                                                                      _T_16959_58 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_15667) begin
                                                                                                                        _T_16959_58 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_15665) begin
                                                                                                                          _T_16959_58 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_15663) begin
                                                                                                                            _T_16959_58 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_15661) begin
                                                                                                                              _T_16959_58 <= _T_9260_58;
                                                                                                                            end else begin
                                                                                                                              _T_16959_58 <= 8'h0;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_58 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_59) begin
        if (_T_15958) begin
          _T_16959_59 <= _T_9260_0;
        end else begin
          if (_T_15956) begin
            _T_16959_59 <= _T_9260_1;
          end else begin
            if (_T_15954) begin
              _T_16959_59 <= _T_9260_2;
            end else begin
              if (_T_15952) begin
                _T_16959_59 <= _T_9260_3;
              end else begin
                if (_T_15950) begin
                  _T_16959_59 <= _T_9260_4;
                end else begin
                  if (_T_15948) begin
                    _T_16959_59 <= _T_9260_5;
                  end else begin
                    if (_T_15946) begin
                      _T_16959_59 <= _T_9260_6;
                    end else begin
                      if (_T_15944) begin
                        _T_16959_59 <= _T_9260_7;
                      end else begin
                        if (_T_15942) begin
                          _T_16959_59 <= _T_9260_8;
                        end else begin
                          if (_T_15940) begin
                            _T_16959_59 <= _T_9260_9;
                          end else begin
                            if (_T_15938) begin
                              _T_16959_59 <= _T_9260_10;
                            end else begin
                              if (_T_15936) begin
                                _T_16959_59 <= _T_9260_11;
                              end else begin
                                if (_T_15934) begin
                                  _T_16959_59 <= _T_9260_12;
                                end else begin
                                  if (_T_15932) begin
                                    _T_16959_59 <= _T_9260_13;
                                  end else begin
                                    if (_T_15930) begin
                                      _T_16959_59 <= _T_9260_14;
                                    end else begin
                                      if (_T_15928) begin
                                        _T_16959_59 <= _T_9260_15;
                                      end else begin
                                        if (_T_15926) begin
                                          _T_16959_59 <= _T_9260_16;
                                        end else begin
                                          if (_T_15924) begin
                                            _T_16959_59 <= _T_9260_17;
                                          end else begin
                                            if (_T_15922) begin
                                              _T_16959_59 <= _T_9260_18;
                                            end else begin
                                              if (_T_15920) begin
                                                _T_16959_59 <= _T_9260_19;
                                              end else begin
                                                if (_T_15918) begin
                                                  _T_16959_59 <= _T_9260_20;
                                                end else begin
                                                  if (_T_15916) begin
                                                    _T_16959_59 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_15914) begin
                                                      _T_16959_59 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_15912) begin
                                                        _T_16959_59 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_15910) begin
                                                          _T_16959_59 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_15908) begin
                                                            _T_16959_59 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_15906) begin
                                                              _T_16959_59 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_15904) begin
                                                                _T_16959_59 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_15902) begin
                                                                  _T_16959_59 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_15900) begin
                                                                    _T_16959_59 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_15898) begin
                                                                      _T_16959_59 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_15896) begin
                                                                        _T_16959_59 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_15894) begin
                                                                          _T_16959_59 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_15892) begin
                                                                            _T_16959_59 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_15890) begin
                                                                              _T_16959_59 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_15888) begin
                                                                                _T_16959_59 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_15886) begin
                                                                                  _T_16959_59 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_15884) begin
                                                                                    _T_16959_59 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_15882) begin
                                                                                      _T_16959_59 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_15880) begin
                                                                                        _T_16959_59 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_15878) begin
                                                                                          _T_16959_59 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_15876) begin
                                                                                            _T_16959_59 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_15874) begin
                                                                                              _T_16959_59 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_15872) begin
                                                                                                _T_16959_59 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_15870) begin
                                                                                                  _T_16959_59 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_15868) begin
                                                                                                    _T_16959_59 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_15866) begin
                                                                                                      _T_16959_59 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_15864) begin
                                                                                                        _T_16959_59 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_15862) begin
                                                                                                          _T_16959_59 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_15860) begin
                                                                                                            _T_16959_59 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_15858) begin
                                                                                                              _T_16959_59 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_15856) begin
                                                                                                                _T_16959_59 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_15854) begin
                                                                                                                  _T_16959_59 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15852) begin
                                                                                                                    _T_16959_59 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_15850) begin
                                                                                                                      _T_16959_59 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_15848) begin
                                                                                                                        _T_16959_59 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_15846) begin
                                                                                                                          _T_16959_59 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_15844) begin
                                                                                                                            _T_16959_59 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_15842) begin
                                                                                                                              _T_16959_59 <= _T_9260_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_15840) begin
                                                                                                                                _T_16959_59 <= _T_9260_59;
                                                                                                                              end else begin
                                                                                                                                _T_16959_59 <= 8'h0;
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_59 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_60) begin
        if (_T_16142) begin
          _T_16959_60 <= _T_9260_0;
        end else begin
          if (_T_16140) begin
            _T_16959_60 <= _T_9260_1;
          end else begin
            if (_T_16138) begin
              _T_16959_60 <= _T_9260_2;
            end else begin
              if (_T_16136) begin
                _T_16959_60 <= _T_9260_3;
              end else begin
                if (_T_16134) begin
                  _T_16959_60 <= _T_9260_4;
                end else begin
                  if (_T_16132) begin
                    _T_16959_60 <= _T_9260_5;
                  end else begin
                    if (_T_16130) begin
                      _T_16959_60 <= _T_9260_6;
                    end else begin
                      if (_T_16128) begin
                        _T_16959_60 <= _T_9260_7;
                      end else begin
                        if (_T_16126) begin
                          _T_16959_60 <= _T_9260_8;
                        end else begin
                          if (_T_16124) begin
                            _T_16959_60 <= _T_9260_9;
                          end else begin
                            if (_T_16122) begin
                              _T_16959_60 <= _T_9260_10;
                            end else begin
                              if (_T_16120) begin
                                _T_16959_60 <= _T_9260_11;
                              end else begin
                                if (_T_16118) begin
                                  _T_16959_60 <= _T_9260_12;
                                end else begin
                                  if (_T_16116) begin
                                    _T_16959_60 <= _T_9260_13;
                                  end else begin
                                    if (_T_16114) begin
                                      _T_16959_60 <= _T_9260_14;
                                    end else begin
                                      if (_T_16112) begin
                                        _T_16959_60 <= _T_9260_15;
                                      end else begin
                                        if (_T_16110) begin
                                          _T_16959_60 <= _T_9260_16;
                                        end else begin
                                          if (_T_16108) begin
                                            _T_16959_60 <= _T_9260_17;
                                          end else begin
                                            if (_T_16106) begin
                                              _T_16959_60 <= _T_9260_18;
                                            end else begin
                                              if (_T_16104) begin
                                                _T_16959_60 <= _T_9260_19;
                                              end else begin
                                                if (_T_16102) begin
                                                  _T_16959_60 <= _T_9260_20;
                                                end else begin
                                                  if (_T_16100) begin
                                                    _T_16959_60 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_16098) begin
                                                      _T_16959_60 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_16096) begin
                                                        _T_16959_60 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_16094) begin
                                                          _T_16959_60 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_16092) begin
                                                            _T_16959_60 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_16090) begin
                                                              _T_16959_60 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_16088) begin
                                                                _T_16959_60 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_16086) begin
                                                                  _T_16959_60 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_16084) begin
                                                                    _T_16959_60 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_16082) begin
                                                                      _T_16959_60 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_16080) begin
                                                                        _T_16959_60 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_16078) begin
                                                                          _T_16959_60 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_16076) begin
                                                                            _T_16959_60 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_16074) begin
                                                                              _T_16959_60 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_16072) begin
                                                                                _T_16959_60 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_16070) begin
                                                                                  _T_16959_60 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_16068) begin
                                                                                    _T_16959_60 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_16066) begin
                                                                                      _T_16959_60 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_16064) begin
                                                                                        _T_16959_60 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_16062) begin
                                                                                          _T_16959_60 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_16060) begin
                                                                                            _T_16959_60 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_16058) begin
                                                                                              _T_16959_60 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_16056) begin
                                                                                                _T_16959_60 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_16054) begin
                                                                                                  _T_16959_60 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_16052) begin
                                                                                                    _T_16959_60 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_16050) begin
                                                                                                      _T_16959_60 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_16048) begin
                                                                                                        _T_16959_60 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_16046) begin
                                                                                                          _T_16959_60 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_16044) begin
                                                                                                            _T_16959_60 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_16042) begin
                                                                                                              _T_16959_60 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_16040) begin
                                                                                                                _T_16959_60 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_16038) begin
                                                                                                                  _T_16959_60 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16036) begin
                                                                                                                    _T_16959_60 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16034) begin
                                                                                                                      _T_16959_60 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16032) begin
                                                                                                                        _T_16959_60 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16030) begin
                                                                                                                          _T_16959_60 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16028) begin
                                                                                                                            _T_16959_60 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16026) begin
                                                                                                                              _T_16959_60 <= _T_9260_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_16024) begin
                                                                                                                                _T_16959_60 <= _T_9260_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_16022) begin
                                                                                                                                  _T_16959_60 <= _T_9260_60;
                                                                                                                                end else begin
                                                                                                                                  _T_16959_60 <= 8'h0;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_60 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_61) begin
        if (_T_16329) begin
          _T_16959_61 <= _T_9260_0;
        end else begin
          if (_T_16327) begin
            _T_16959_61 <= _T_9260_1;
          end else begin
            if (_T_16325) begin
              _T_16959_61 <= _T_9260_2;
            end else begin
              if (_T_16323) begin
                _T_16959_61 <= _T_9260_3;
              end else begin
                if (_T_16321) begin
                  _T_16959_61 <= _T_9260_4;
                end else begin
                  if (_T_16319) begin
                    _T_16959_61 <= _T_9260_5;
                  end else begin
                    if (_T_16317) begin
                      _T_16959_61 <= _T_9260_6;
                    end else begin
                      if (_T_16315) begin
                        _T_16959_61 <= _T_9260_7;
                      end else begin
                        if (_T_16313) begin
                          _T_16959_61 <= _T_9260_8;
                        end else begin
                          if (_T_16311) begin
                            _T_16959_61 <= _T_9260_9;
                          end else begin
                            if (_T_16309) begin
                              _T_16959_61 <= _T_9260_10;
                            end else begin
                              if (_T_16307) begin
                                _T_16959_61 <= _T_9260_11;
                              end else begin
                                if (_T_16305) begin
                                  _T_16959_61 <= _T_9260_12;
                                end else begin
                                  if (_T_16303) begin
                                    _T_16959_61 <= _T_9260_13;
                                  end else begin
                                    if (_T_16301) begin
                                      _T_16959_61 <= _T_9260_14;
                                    end else begin
                                      if (_T_16299) begin
                                        _T_16959_61 <= _T_9260_15;
                                      end else begin
                                        if (_T_16297) begin
                                          _T_16959_61 <= _T_9260_16;
                                        end else begin
                                          if (_T_16295) begin
                                            _T_16959_61 <= _T_9260_17;
                                          end else begin
                                            if (_T_16293) begin
                                              _T_16959_61 <= _T_9260_18;
                                            end else begin
                                              if (_T_16291) begin
                                                _T_16959_61 <= _T_9260_19;
                                              end else begin
                                                if (_T_16289) begin
                                                  _T_16959_61 <= _T_9260_20;
                                                end else begin
                                                  if (_T_16287) begin
                                                    _T_16959_61 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_16285) begin
                                                      _T_16959_61 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_16283) begin
                                                        _T_16959_61 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_16281) begin
                                                          _T_16959_61 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_16279) begin
                                                            _T_16959_61 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_16277) begin
                                                              _T_16959_61 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_16275) begin
                                                                _T_16959_61 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_16273) begin
                                                                  _T_16959_61 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_16271) begin
                                                                    _T_16959_61 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_16269) begin
                                                                      _T_16959_61 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_16267) begin
                                                                        _T_16959_61 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_16265) begin
                                                                          _T_16959_61 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_16263) begin
                                                                            _T_16959_61 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_16261) begin
                                                                              _T_16959_61 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_16259) begin
                                                                                _T_16959_61 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_16257) begin
                                                                                  _T_16959_61 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_16255) begin
                                                                                    _T_16959_61 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_16253) begin
                                                                                      _T_16959_61 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_16251) begin
                                                                                        _T_16959_61 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_16249) begin
                                                                                          _T_16959_61 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_16247) begin
                                                                                            _T_16959_61 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_16245) begin
                                                                                              _T_16959_61 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_16243) begin
                                                                                                _T_16959_61 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_16241) begin
                                                                                                  _T_16959_61 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_16239) begin
                                                                                                    _T_16959_61 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_16237) begin
                                                                                                      _T_16959_61 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_16235) begin
                                                                                                        _T_16959_61 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_16233) begin
                                                                                                          _T_16959_61 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_16231) begin
                                                                                                            _T_16959_61 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_16229) begin
                                                                                                              _T_16959_61 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_16227) begin
                                                                                                                _T_16959_61 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_16225) begin
                                                                                                                  _T_16959_61 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16223) begin
                                                                                                                    _T_16959_61 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16221) begin
                                                                                                                      _T_16959_61 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16219) begin
                                                                                                                        _T_16959_61 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16217) begin
                                                                                                                          _T_16959_61 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16215) begin
                                                                                                                            _T_16959_61 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16213) begin
                                                                                                                              _T_16959_61 <= _T_9260_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_16211) begin
                                                                                                                                _T_16959_61 <= _T_9260_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_16209) begin
                                                                                                                                  _T_16959_61 <= _T_9260_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_16207) begin
                                                                                                                                    _T_16959_61 <= _T_9260_61;
                                                                                                                                  end else begin
                                                                                                                                    _T_16959_61 <= 8'h0;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_61 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_62) begin
        if (_T_16519) begin
          _T_16959_62 <= _T_9260_0;
        end else begin
          if (_T_16517) begin
            _T_16959_62 <= _T_9260_1;
          end else begin
            if (_T_16515) begin
              _T_16959_62 <= _T_9260_2;
            end else begin
              if (_T_16513) begin
                _T_16959_62 <= _T_9260_3;
              end else begin
                if (_T_16511) begin
                  _T_16959_62 <= _T_9260_4;
                end else begin
                  if (_T_16509) begin
                    _T_16959_62 <= _T_9260_5;
                  end else begin
                    if (_T_16507) begin
                      _T_16959_62 <= _T_9260_6;
                    end else begin
                      if (_T_16505) begin
                        _T_16959_62 <= _T_9260_7;
                      end else begin
                        if (_T_16503) begin
                          _T_16959_62 <= _T_9260_8;
                        end else begin
                          if (_T_16501) begin
                            _T_16959_62 <= _T_9260_9;
                          end else begin
                            if (_T_16499) begin
                              _T_16959_62 <= _T_9260_10;
                            end else begin
                              if (_T_16497) begin
                                _T_16959_62 <= _T_9260_11;
                              end else begin
                                if (_T_16495) begin
                                  _T_16959_62 <= _T_9260_12;
                                end else begin
                                  if (_T_16493) begin
                                    _T_16959_62 <= _T_9260_13;
                                  end else begin
                                    if (_T_16491) begin
                                      _T_16959_62 <= _T_9260_14;
                                    end else begin
                                      if (_T_16489) begin
                                        _T_16959_62 <= _T_9260_15;
                                      end else begin
                                        if (_T_16487) begin
                                          _T_16959_62 <= _T_9260_16;
                                        end else begin
                                          if (_T_16485) begin
                                            _T_16959_62 <= _T_9260_17;
                                          end else begin
                                            if (_T_16483) begin
                                              _T_16959_62 <= _T_9260_18;
                                            end else begin
                                              if (_T_16481) begin
                                                _T_16959_62 <= _T_9260_19;
                                              end else begin
                                                if (_T_16479) begin
                                                  _T_16959_62 <= _T_9260_20;
                                                end else begin
                                                  if (_T_16477) begin
                                                    _T_16959_62 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_16475) begin
                                                      _T_16959_62 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_16473) begin
                                                        _T_16959_62 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_16471) begin
                                                          _T_16959_62 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_16469) begin
                                                            _T_16959_62 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_16467) begin
                                                              _T_16959_62 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_16465) begin
                                                                _T_16959_62 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_16463) begin
                                                                  _T_16959_62 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_16461) begin
                                                                    _T_16959_62 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_16459) begin
                                                                      _T_16959_62 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_16457) begin
                                                                        _T_16959_62 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_16455) begin
                                                                          _T_16959_62 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_16453) begin
                                                                            _T_16959_62 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_16451) begin
                                                                              _T_16959_62 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_16449) begin
                                                                                _T_16959_62 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_16447) begin
                                                                                  _T_16959_62 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_16445) begin
                                                                                    _T_16959_62 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_16443) begin
                                                                                      _T_16959_62 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_16441) begin
                                                                                        _T_16959_62 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_16439) begin
                                                                                          _T_16959_62 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_16437) begin
                                                                                            _T_16959_62 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_16435) begin
                                                                                              _T_16959_62 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_16433) begin
                                                                                                _T_16959_62 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_16431) begin
                                                                                                  _T_16959_62 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_16429) begin
                                                                                                    _T_16959_62 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_16427) begin
                                                                                                      _T_16959_62 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_16425) begin
                                                                                                        _T_16959_62 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_16423) begin
                                                                                                          _T_16959_62 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_16421) begin
                                                                                                            _T_16959_62 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_16419) begin
                                                                                                              _T_16959_62 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_16417) begin
                                                                                                                _T_16959_62 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_16415) begin
                                                                                                                  _T_16959_62 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16413) begin
                                                                                                                    _T_16959_62 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16411) begin
                                                                                                                      _T_16959_62 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16409) begin
                                                                                                                        _T_16959_62 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16407) begin
                                                                                                                          _T_16959_62 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16405) begin
                                                                                                                            _T_16959_62 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16403) begin
                                                                                                                              _T_16959_62 <= _T_9260_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_16401) begin
                                                                                                                                _T_16959_62 <= _T_9260_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_16399) begin
                                                                                                                                  _T_16959_62 <= _T_9260_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_16397) begin
                                                                                                                                    _T_16959_62 <= _T_9260_61;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_16395) begin
                                                                                                                                      _T_16959_62 <= _T_9260_62;
                                                                                                                                    end else begin
                                                                                                                                      _T_16959_62 <= 8'h0;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_62 <= 8'h0;
      end
    end
    if (_T_9256) begin
      if (_T_9330_63) begin
        if (_T_16712) begin
          _T_16959_63 <= _T_9260_0;
        end else begin
          if (_T_16710) begin
            _T_16959_63 <= _T_9260_1;
          end else begin
            if (_T_16708) begin
              _T_16959_63 <= _T_9260_2;
            end else begin
              if (_T_16706) begin
                _T_16959_63 <= _T_9260_3;
              end else begin
                if (_T_16704) begin
                  _T_16959_63 <= _T_9260_4;
                end else begin
                  if (_T_16702) begin
                    _T_16959_63 <= _T_9260_5;
                  end else begin
                    if (_T_16700) begin
                      _T_16959_63 <= _T_9260_6;
                    end else begin
                      if (_T_16698) begin
                        _T_16959_63 <= _T_9260_7;
                      end else begin
                        if (_T_16696) begin
                          _T_16959_63 <= _T_9260_8;
                        end else begin
                          if (_T_16694) begin
                            _T_16959_63 <= _T_9260_9;
                          end else begin
                            if (_T_16692) begin
                              _T_16959_63 <= _T_9260_10;
                            end else begin
                              if (_T_16690) begin
                                _T_16959_63 <= _T_9260_11;
                              end else begin
                                if (_T_16688) begin
                                  _T_16959_63 <= _T_9260_12;
                                end else begin
                                  if (_T_16686) begin
                                    _T_16959_63 <= _T_9260_13;
                                  end else begin
                                    if (_T_16684) begin
                                      _T_16959_63 <= _T_9260_14;
                                    end else begin
                                      if (_T_16682) begin
                                        _T_16959_63 <= _T_9260_15;
                                      end else begin
                                        if (_T_16680) begin
                                          _T_16959_63 <= _T_9260_16;
                                        end else begin
                                          if (_T_16678) begin
                                            _T_16959_63 <= _T_9260_17;
                                          end else begin
                                            if (_T_16676) begin
                                              _T_16959_63 <= _T_9260_18;
                                            end else begin
                                              if (_T_16674) begin
                                                _T_16959_63 <= _T_9260_19;
                                              end else begin
                                                if (_T_16672) begin
                                                  _T_16959_63 <= _T_9260_20;
                                                end else begin
                                                  if (_T_16670) begin
                                                    _T_16959_63 <= _T_9260_21;
                                                  end else begin
                                                    if (_T_16668) begin
                                                      _T_16959_63 <= _T_9260_22;
                                                    end else begin
                                                      if (_T_16666) begin
                                                        _T_16959_63 <= _T_9260_23;
                                                      end else begin
                                                        if (_T_16664) begin
                                                          _T_16959_63 <= _T_9260_24;
                                                        end else begin
                                                          if (_T_16662) begin
                                                            _T_16959_63 <= _T_9260_25;
                                                          end else begin
                                                            if (_T_16660) begin
                                                              _T_16959_63 <= _T_9260_26;
                                                            end else begin
                                                              if (_T_16658) begin
                                                                _T_16959_63 <= _T_9260_27;
                                                              end else begin
                                                                if (_T_16656) begin
                                                                  _T_16959_63 <= _T_9260_28;
                                                                end else begin
                                                                  if (_T_16654) begin
                                                                    _T_16959_63 <= _T_9260_29;
                                                                  end else begin
                                                                    if (_T_16652) begin
                                                                      _T_16959_63 <= _T_9260_30;
                                                                    end else begin
                                                                      if (_T_16650) begin
                                                                        _T_16959_63 <= _T_9260_31;
                                                                      end else begin
                                                                        if (_T_16648) begin
                                                                          _T_16959_63 <= _T_9260_32;
                                                                        end else begin
                                                                          if (_T_16646) begin
                                                                            _T_16959_63 <= _T_9260_33;
                                                                          end else begin
                                                                            if (_T_16644) begin
                                                                              _T_16959_63 <= _T_9260_34;
                                                                            end else begin
                                                                              if (_T_16642) begin
                                                                                _T_16959_63 <= _T_9260_35;
                                                                              end else begin
                                                                                if (_T_16640) begin
                                                                                  _T_16959_63 <= _T_9260_36;
                                                                                end else begin
                                                                                  if (_T_16638) begin
                                                                                    _T_16959_63 <= _T_9260_37;
                                                                                  end else begin
                                                                                    if (_T_16636) begin
                                                                                      _T_16959_63 <= _T_9260_38;
                                                                                    end else begin
                                                                                      if (_T_16634) begin
                                                                                        _T_16959_63 <= _T_9260_39;
                                                                                      end else begin
                                                                                        if (_T_16632) begin
                                                                                          _T_16959_63 <= _T_9260_40;
                                                                                        end else begin
                                                                                          if (_T_16630) begin
                                                                                            _T_16959_63 <= _T_9260_41;
                                                                                          end else begin
                                                                                            if (_T_16628) begin
                                                                                              _T_16959_63 <= _T_9260_42;
                                                                                            end else begin
                                                                                              if (_T_16626) begin
                                                                                                _T_16959_63 <= _T_9260_43;
                                                                                              end else begin
                                                                                                if (_T_16624) begin
                                                                                                  _T_16959_63 <= _T_9260_44;
                                                                                                end else begin
                                                                                                  if (_T_16622) begin
                                                                                                    _T_16959_63 <= _T_9260_45;
                                                                                                  end else begin
                                                                                                    if (_T_16620) begin
                                                                                                      _T_16959_63 <= _T_9260_46;
                                                                                                    end else begin
                                                                                                      if (_T_16618) begin
                                                                                                        _T_16959_63 <= _T_9260_47;
                                                                                                      end else begin
                                                                                                        if (_T_16616) begin
                                                                                                          _T_16959_63 <= _T_9260_48;
                                                                                                        end else begin
                                                                                                          if (_T_16614) begin
                                                                                                            _T_16959_63 <= _T_9260_49;
                                                                                                          end else begin
                                                                                                            if (_T_16612) begin
                                                                                                              _T_16959_63 <= _T_9260_50;
                                                                                                            end else begin
                                                                                                              if (_T_16610) begin
                                                                                                                _T_16959_63 <= _T_9260_51;
                                                                                                              end else begin
                                                                                                                if (_T_16608) begin
                                                                                                                  _T_16959_63 <= _T_9260_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16606) begin
                                                                                                                    _T_16959_63 <= _T_9260_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16604) begin
                                                                                                                      _T_16959_63 <= _T_9260_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16602) begin
                                                                                                                        _T_16959_63 <= _T_9260_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16600) begin
                                                                                                                          _T_16959_63 <= _T_9260_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16598) begin
                                                                                                                            _T_16959_63 <= _T_9260_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16596) begin
                                                                                                                              _T_16959_63 <= _T_9260_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_16594) begin
                                                                                                                                _T_16959_63 <= _T_9260_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_16592) begin
                                                                                                                                  _T_16959_63 <= _T_9260_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_16590) begin
                                                                                                                                    _T_16959_63 <= _T_9260_61;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_16588) begin
                                                                                                                                      _T_16959_63 <= _T_9260_62;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_16586) begin
                                                                                                                                        _T_16959_63 <= _T_9260_63;
                                                                                                                                      end else begin
                                                                                                                                        _T_16959_63 <= 8'h0;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_16959_63 <= 8'h0;
      end
    end
    if (_T_326) begin
      _T_17290 <= 1'h0;
    end else begin
      _T_17290 <= _T_16716;
    end
    if (_T_16716) begin
      _T_17294_0 <= _T_17161;
    end
    if (_T_16716) begin
      _T_17294_1 <= _T_17163;
    end
    if (_T_16716) begin
      _T_17294_2 <= _T_17165;
    end
    if (_T_16716) begin
      _T_17294_3 <= _T_17167;
    end
    if (_T_16716) begin
      _T_17294_4 <= _T_17169;
    end
    if (_T_16716) begin
      _T_17294_5 <= _T_17171;
    end
    if (_T_16716) begin
      _T_17294_6 <= _T_17173;
    end
    if (_T_16716) begin
      _T_17294_7 <= _T_17175;
    end
    if (_T_16716) begin
      _T_17294_8 <= _T_17177;
    end
    if (_T_16716) begin
      _T_17294_9 <= _T_17179;
    end
    if (_T_16716) begin
      _T_17294_10 <= _T_17181;
    end
    if (_T_16716) begin
      _T_17294_11 <= _T_17183;
    end
    if (_T_16716) begin
      _T_17294_12 <= _T_17185;
    end
    if (_T_16716) begin
      _T_17294_13 <= _T_17187;
    end
    if (_T_16716) begin
      _T_17294_14 <= _T_17189;
    end
    if (_T_16716) begin
      _T_17294_15 <= _T_17191;
    end
    if (_T_16716) begin
      _T_17294_16 <= _T_17193;
    end
    if (_T_16716) begin
      _T_17294_17 <= _T_17195;
    end
    if (_T_16716) begin
      _T_17294_18 <= _T_17197;
    end
    if (_T_16716) begin
      _T_17294_19 <= _T_17199;
    end
    if (_T_16716) begin
      _T_17294_20 <= _T_17201;
    end
    if (_T_16716) begin
      _T_17294_21 <= _T_17203;
    end
    if (_T_16716) begin
      _T_17294_22 <= _T_17205;
    end
    if (_T_16716) begin
      _T_17294_23 <= _T_17207;
    end
    if (_T_16716) begin
      _T_17294_24 <= _T_17209;
    end
    if (_T_16716) begin
      _T_17294_25 <= _T_17211;
    end
    if (_T_16716) begin
      _T_17294_26 <= _T_17213;
    end
    if (_T_16716) begin
      _T_17294_27 <= _T_17215;
    end
    if (_T_16716) begin
      _T_17294_28 <= _T_17217;
    end
    if (_T_16716) begin
      _T_17294_29 <= _T_17219;
    end
    if (_T_16716) begin
      _T_17294_30 <= _T_17221;
    end
    if (_T_16716) begin
      _T_17294_31 <= _T_17223;
    end
    if (_T_16716) begin
      _T_17294_32 <= _T_17225;
    end
    if (_T_16716) begin
      _T_17294_33 <= _T_17227;
    end
    if (_T_16716) begin
      _T_17294_34 <= _T_17229;
    end
    if (_T_16716) begin
      _T_17294_35 <= _T_17231;
    end
    if (_T_16716) begin
      _T_17294_36 <= _T_17233;
    end
    if (_T_16716) begin
      _T_17294_37 <= _T_17235;
    end
    if (_T_16716) begin
      _T_17294_38 <= _T_17237;
    end
    if (_T_16716) begin
      _T_17294_39 <= _T_17239;
    end
    if (_T_16716) begin
      _T_17294_40 <= _T_17241;
    end
    if (_T_16716) begin
      _T_17294_41 <= _T_17243;
    end
    if (_T_16716) begin
      _T_17294_42 <= _T_17245;
    end
    if (_T_16716) begin
      _T_17294_43 <= _T_17247;
    end
    if (_T_16716) begin
      _T_17294_44 <= _T_17249;
    end
    if (_T_16716) begin
      _T_17294_45 <= _T_17251;
    end
    if (_T_16716) begin
      _T_17294_46 <= _T_17253;
    end
    if (_T_16716) begin
      _T_17294_47 <= _T_17255;
    end
    if (_T_16716) begin
      _T_17294_48 <= _T_17257;
    end
    if (_T_16716) begin
      _T_17294_49 <= _T_17259;
    end
    if (_T_16716) begin
      _T_17294_50 <= _T_17261;
    end
    if (_T_16716) begin
      _T_17294_51 <= _T_17263;
    end
    if (_T_16716) begin
      _T_17294_52 <= _T_17265;
    end
    if (_T_16716) begin
      _T_17294_53 <= _T_17267;
    end
    if (_T_16716) begin
      _T_17294_54 <= _T_17269;
    end
    if (_T_16716) begin
      _T_17294_55 <= _T_17271;
    end
    if (_T_16716) begin
      _T_17294_56 <= _T_17273;
    end
    if (_T_16716) begin
      _T_17294_57 <= _T_17275;
    end
    if (_T_16716) begin
      _T_17294_58 <= _T_17277;
    end
    if (_T_16716) begin
      _T_17294_59 <= _T_17279;
    end
    if (_T_16716) begin
      _T_17294_60 <= _T_17281;
    end
    if (_T_16716) begin
      _T_17294_61 <= _T_17283;
    end
    if (_T_16716) begin
      _T_17294_62 <= _T_17285;
    end
    if (_T_16716) begin
      _T_17294_63 <= _T_17287;
    end
    if (_T_326) begin
      _T_17499_0 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_0 <= _T_16855_0;
      end
    end
    if (_T_326) begin
      _T_17499_1 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_1 <= _T_16855_1;
      end
    end
    if (_T_326) begin
      _T_17499_2 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_2 <= _T_16855_2;
      end
    end
    if (_T_326) begin
      _T_17499_3 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_3 <= _T_16855_3;
      end
    end
    if (_T_326) begin
      _T_17499_4 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_4 <= _T_16855_4;
      end
    end
    if (_T_326) begin
      _T_17499_5 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_5 <= _T_16855_5;
      end
    end
    if (_T_326) begin
      _T_17499_6 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_6 <= _T_16855_6;
      end
    end
    if (_T_326) begin
      _T_17499_7 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_7 <= _T_16855_7;
      end
    end
    if (_T_326) begin
      _T_17499_8 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_8 <= _T_16855_8;
      end
    end
    if (_T_326) begin
      _T_17499_9 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_9 <= _T_16855_9;
      end
    end
    if (_T_326) begin
      _T_17499_10 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_10 <= _T_16855_10;
      end
    end
    if (_T_326) begin
      _T_17499_11 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_11 <= _T_16855_11;
      end
    end
    if (_T_326) begin
      _T_17499_12 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_12 <= _T_16855_12;
      end
    end
    if (_T_326) begin
      _T_17499_13 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_13 <= _T_16855_13;
      end
    end
    if (_T_326) begin
      _T_17499_14 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_14 <= _T_16855_14;
      end
    end
    if (_T_326) begin
      _T_17499_15 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_15 <= _T_16855_15;
      end
    end
    if (_T_326) begin
      _T_17499_16 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_16 <= _T_16855_16;
      end
    end
    if (_T_326) begin
      _T_17499_17 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_17 <= _T_16855_17;
      end
    end
    if (_T_326) begin
      _T_17499_18 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_18 <= _T_16855_18;
      end
    end
    if (_T_326) begin
      _T_17499_19 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_19 <= _T_16855_19;
      end
    end
    if (_T_326) begin
      _T_17499_20 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_20 <= _T_16855_20;
      end
    end
    if (_T_326) begin
      _T_17499_21 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_21 <= _T_16855_21;
      end
    end
    if (_T_326) begin
      _T_17499_22 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_22 <= _T_16855_22;
      end
    end
    if (_T_326) begin
      _T_17499_23 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_23 <= _T_16855_23;
      end
    end
    if (_T_326) begin
      _T_17499_24 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_24 <= _T_16855_24;
      end
    end
    if (_T_326) begin
      _T_17499_25 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_25 <= _T_16855_25;
      end
    end
    if (_T_326) begin
      _T_17499_26 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_26 <= _T_16855_26;
      end
    end
    if (_T_326) begin
      _T_17499_27 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_27 <= _T_16855_27;
      end
    end
    if (_T_326) begin
      _T_17499_28 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_28 <= _T_16855_28;
      end
    end
    if (_T_326) begin
      _T_17499_29 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_29 <= _T_16855_29;
      end
    end
    if (_T_326) begin
      _T_17499_30 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_30 <= _T_16855_30;
      end
    end
    if (_T_326) begin
      _T_17499_31 <= 1'h0;
    end else begin
      if (_T_16716) begin
        _T_17499_31 <= _T_16855_31;
      end
    end
    if (_T_16716) begin
      _T_17603_0 <= _T_16959_0;
    end
    if (_T_16716) begin
      _T_17603_1 <= _T_16959_1;
    end
    if (_T_16716) begin
      _T_17603_2 <= _T_16959_2;
    end
    if (_T_16716) begin
      _T_17603_3 <= _T_16959_3;
    end
    if (_T_16716) begin
      _T_17603_4 <= _T_16959_4;
    end
    if (_T_16716) begin
      _T_17603_5 <= _T_16959_5;
    end
    if (_T_16716) begin
      _T_17603_6 <= _T_16959_6;
    end
    if (_T_16716) begin
      _T_17603_7 <= _T_16959_7;
    end
    if (_T_16716) begin
      _T_17603_8 <= _T_16959_8;
    end
    if (_T_16716) begin
      _T_17603_9 <= _T_16959_9;
    end
    if (_T_16716) begin
      _T_17603_10 <= _T_16959_10;
    end
    if (_T_16716) begin
      _T_17603_11 <= _T_16959_11;
    end
    if (_T_16716) begin
      _T_17603_12 <= _T_16959_12;
    end
    if (_T_16716) begin
      _T_17603_13 <= _T_16959_13;
    end
    if (_T_16716) begin
      _T_17603_14 <= _T_16959_14;
    end
    if (_T_16716) begin
      _T_17603_15 <= _T_16959_15;
    end
    if (_T_16716) begin
      _T_17603_16 <= _T_16959_16;
    end
    if (_T_16716) begin
      _T_17603_17 <= _T_16959_17;
    end
    if (_T_16716) begin
      _T_17603_18 <= _T_16959_18;
    end
    if (_T_16716) begin
      _T_17603_19 <= _T_16959_19;
    end
    if (_T_16716) begin
      _T_17603_20 <= _T_16959_20;
    end
    if (_T_16716) begin
      _T_17603_21 <= _T_16959_21;
    end
    if (_T_16716) begin
      _T_17603_22 <= _T_16959_22;
    end
    if (_T_16716) begin
      _T_17603_23 <= _T_16959_23;
    end
    if (_T_16716) begin
      _T_17603_24 <= _T_16959_24;
    end
    if (_T_16716) begin
      _T_17603_25 <= _T_16959_25;
    end
    if (_T_16716) begin
      _T_17603_26 <= _T_16959_26;
    end
    if (_T_16716) begin
      _T_17603_27 <= _T_16959_27;
    end
    if (_T_16716) begin
      _T_17603_28 <= _T_16959_28;
    end
    if (_T_16716) begin
      _T_17603_29 <= _T_16959_29;
    end
    if (_T_16716) begin
      _T_17603_30 <= _T_16959_30;
    end
    if (_T_16716) begin
      _T_17603_31 <= _T_16959_31;
    end
    if (_T_16716) begin
      _T_17603_32 <= _T_16959_32;
    end
    if (_T_16716) begin
      _T_17603_33 <= _T_16959_33;
    end
    if (_T_16716) begin
      _T_17603_34 <= _T_16959_34;
    end
    if (_T_16716) begin
      _T_17603_35 <= _T_16959_35;
    end
    if (_T_16716) begin
      _T_17603_36 <= _T_16959_36;
    end
    if (_T_16716) begin
      _T_17603_37 <= _T_16959_37;
    end
    if (_T_16716) begin
      _T_17603_38 <= _T_16959_38;
    end
    if (_T_16716) begin
      _T_17603_39 <= _T_16959_39;
    end
    if (_T_16716) begin
      _T_17603_40 <= _T_16959_40;
    end
    if (_T_16716) begin
      _T_17603_41 <= _T_16959_41;
    end
    if (_T_16716) begin
      _T_17603_42 <= _T_16959_42;
    end
    if (_T_16716) begin
      _T_17603_43 <= _T_16959_43;
    end
    if (_T_16716) begin
      _T_17603_44 <= _T_16959_44;
    end
    if (_T_16716) begin
      _T_17603_45 <= _T_16959_45;
    end
    if (_T_16716) begin
      _T_17603_46 <= _T_16959_46;
    end
    if (_T_16716) begin
      _T_17603_47 <= _T_16959_47;
    end
    if (_T_16716) begin
      _T_17603_48 <= _T_16959_48;
    end
    if (_T_16716) begin
      _T_17603_49 <= _T_16959_49;
    end
    if (_T_16716) begin
      _T_17603_50 <= _T_16959_50;
    end
    if (_T_16716) begin
      _T_17603_51 <= _T_16959_51;
    end
    if (_T_16716) begin
      _T_17603_52 <= _T_16959_52;
    end
    if (_T_16716) begin
      _T_17603_53 <= _T_16959_53;
    end
    if (_T_16716) begin
      _T_17603_54 <= _T_16959_54;
    end
    if (_T_16716) begin
      _T_17603_55 <= _T_16959_55;
    end
    if (_T_16716) begin
      _T_17603_56 <= _T_16959_56;
    end
    if (_T_16716) begin
      _T_17603_57 <= _T_16959_57;
    end
    if (_T_16716) begin
      _T_17603_58 <= _T_16959_58;
    end
    if (_T_16716) begin
      _T_17603_59 <= _T_16959_59;
    end
    if (_T_16716) begin
      _T_17603_60 <= _T_16959_60;
    end
    if (_T_16716) begin
      _T_17603_61 <= _T_16959_61;
    end
    if (_T_16716) begin
      _T_17603_62 <= _T_16959_62;
    end
    if (_T_16716) begin
      _T_17603_63 <= _T_16959_63;
    end
  end
endmodule
